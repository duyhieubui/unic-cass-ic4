magic
tech sky130A
magscale 1 2
timestamp 1698980770
<< metal2 >>
rect 110620 16000 111020 16010
rect 114830 16000 115230 16010
rect 119260 16000 119660 16010
rect 123620 16000 124020 16010
rect 128100 16000 128500 16010
rect 111020 15600 111030 16000
rect 110620 15500 111030 15600
rect 111020 15100 111030 15500
rect 110620 15000 111030 15100
rect 111020 14600 111030 15000
rect 110620 14500 111030 14600
rect 111020 14100 111030 14500
rect 110620 14000 111030 14100
rect 111020 13600 111030 14000
rect 110620 13500 111030 13600
rect 111020 13100 111030 13500
rect 110620 13000 111030 13100
rect 111020 12600 111030 13000
rect 110620 12500 111030 12600
rect 111020 12100 111030 12500
rect 110620 2401 111030 12100
rect 115230 15600 115250 16000
rect 114830 15500 115250 15600
rect 115230 15100 115250 15500
rect 114830 15000 115250 15100
rect 115230 14600 115250 15000
rect 114830 14500 115250 14600
rect 115230 14100 115250 14500
rect 114830 14000 115250 14100
rect 115230 13600 115250 14000
rect 114830 13500 115250 13600
rect 115230 13100 115250 13500
rect 114830 13000 115250 13100
rect 115230 12600 115250 13000
rect 114830 12500 115250 12600
rect 115230 12100 115250 12500
rect 114830 4409 115250 12100
rect 119660 15600 119670 16000
rect 119260 15500 119670 15600
rect 119660 15100 119670 15500
rect 119260 15000 119670 15100
rect 119660 14600 119670 15000
rect 119260 14500 119670 14600
rect 119660 14100 119670 14500
rect 119260 14000 119670 14100
rect 119660 13600 119670 14000
rect 119260 13500 119670 13600
rect 119660 13100 119670 13500
rect 119260 13000 119670 13100
rect 119660 12600 119670 13000
rect 119260 12500 119670 12600
rect 119660 12100 119670 12500
rect 119260 6399 119670 12100
rect 124020 15600 124030 16000
rect 123620 15500 124030 15600
rect 124020 15100 124030 15500
rect 123620 15000 124030 15100
rect 124020 14600 124030 15000
rect 123620 14500 124030 14600
rect 124020 14100 124030 14500
rect 123620 14000 124030 14100
rect 124020 13600 124030 14000
rect 123620 13500 124030 13600
rect 124020 13100 124030 13500
rect 123620 13000 124030 13100
rect 124020 12600 124030 13000
rect 123620 12500 124030 12600
rect 124020 12100 124030 12500
rect 123620 8400 124030 12100
rect 128500 15600 128510 16000
rect 128100 15500 128510 15600
rect 128500 15100 128510 15500
rect 128100 15000 128510 15100
rect 128500 14600 128510 15000
rect 128100 14500 128510 14600
rect 128500 14100 128510 14500
rect 128100 14000 128510 14100
rect 128500 13600 128510 14000
rect 128100 13500 128510 13600
rect 128500 13100 128510 13500
rect 128100 13000 128510 13100
rect 128500 12600 128510 13000
rect 128100 12500 128510 12600
rect 128500 12100 128510 12500
rect 128100 10400 128510 12100
rect 144582 14500 144982 14536
rect 144582 14000 144982 14100
rect 144582 13500 144982 13600
rect 144582 13000 144982 13100
rect 144582 12500 144982 12600
rect 128100 10000 141432 10400
rect 123620 8000 137882 8400
rect 119260 6000 134340 6399
rect 114830 4009 130800 4409
rect 114830 4000 119252 4009
rect 126744 4000 130800 4009
rect 110620 2000 127250 2401
rect 126850 790 127250 2000
rect 126860 780 127250 790
rect 126870 770 127240 780
rect 126880 760 127230 770
rect 126890 750 127220 760
rect 126900 740 127210 750
rect 130390 740 130800 4000
rect 133940 740 134340 6000
rect 137482 740 137882 8000
rect 141032 780 141432 10000
rect 144582 810 144982 12100
rect 144592 800 144982 810
rect 144602 790 144972 800
rect 144612 780 144962 790
rect 141042 770 141432 780
rect 144622 770 144952 780
rect 141052 760 141422 770
rect 144632 760 144942 770
rect 141062 750 141412 760
rect 144642 750 144932 760
rect 141072 740 141402 750
rect 144652 740 144922 750
rect 126910 730 127200 740
rect 130400 730 130800 740
rect 133950 730 134340 740
rect 137492 730 137882 740
rect 141082 730 141392 740
rect 144662 730 144912 740
rect 126920 720 127190 730
rect 130410 720 130790 730
rect 133960 720 134330 730
rect 137502 720 137872 730
rect 141092 720 141382 730
rect 144672 720 144902 730
rect 126930 710 127180 720
rect 130420 710 130780 720
rect 133970 710 134320 720
rect 137512 710 137862 720
rect 141102 710 141372 720
rect 144682 710 144892 720
rect 126940 700 127170 710
rect 130430 700 130770 710
rect 133980 700 134310 710
rect 137522 700 137852 710
rect 141112 700 141362 710
rect 144692 700 144882 710
rect 126950 690 127160 700
rect 130440 690 130760 700
rect 133990 690 134300 700
rect 137532 690 137842 700
rect 141122 690 141352 700
rect 144702 690 144872 700
rect 126960 680 127150 690
rect 130450 680 130750 690
rect 134000 680 134290 690
rect 137542 680 137832 690
rect 141132 680 141342 690
rect 144712 680 144862 690
rect 126970 670 127140 680
rect 130460 670 130740 680
rect 134010 670 134280 680
rect 137552 670 137822 680
rect 141142 670 141332 680
rect 144722 670 144852 680
rect 126980 660 127130 670
rect 130470 660 130730 670
rect 134020 660 134270 670
rect 137562 660 137812 670
rect 141152 660 141322 670
rect 126990 650 127120 660
rect 130480 650 130720 660
rect 134030 650 134260 660
rect 137572 650 137802 660
rect 141162 650 141312 660
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 650
rect 130490 640 130710 650
rect 134040 640 134250 650
rect 137582 640 137792 650
rect 141172 640 141302 650
rect 130500 630 130700 640
rect 134050 630 134240 640
rect 137592 630 137782 640
rect 130510 620 130690 630
rect 134060 620 134230 630
rect 137602 620 137772 630
rect 130520 610 130680 620
rect 134070 610 134220 620
rect 137612 610 137762 620
rect 130530 600 130670 610
rect 134080 600 134210 610
rect 137622 600 137752 610
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 600
rect 131726 -800 131838 480
rect 132908 -800 133020 600
rect 134090 -800 134202 600
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 600
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 640
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 670
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 110620 15600 111020 16000
rect 110620 15100 111020 15500
rect 110620 14600 111020 15000
rect 110620 14100 111020 14500
rect 110620 13600 111020 14000
rect 110620 13100 111020 13500
rect 110620 12600 111020 13000
rect 110620 12100 111020 12500
rect 114830 15600 115230 16000
rect 114830 15100 115230 15500
rect 114830 14600 115230 15000
rect 114830 14100 115230 14500
rect 114830 13600 115230 14000
rect 114830 13100 115230 13500
rect 114830 12600 115230 13000
rect 114830 12100 115230 12500
rect 119260 15600 119660 16000
rect 119260 15100 119660 15500
rect 119260 14600 119660 15000
rect 119260 14100 119660 14500
rect 119260 13600 119660 14000
rect 119260 13100 119660 13500
rect 119260 12600 119660 13000
rect 119260 12100 119660 12500
rect 123620 15600 124020 16000
rect 123620 15100 124020 15500
rect 123620 14600 124020 15000
rect 123620 14100 124020 14500
rect 123620 13600 124020 14000
rect 123620 13100 124020 13500
rect 123620 12600 124020 13000
rect 123620 12100 124020 12500
rect 128100 15600 128500 16000
rect 128100 15100 128500 15500
rect 128100 14600 128500 15000
rect 128100 14100 128500 14500
rect 128100 13600 128500 14000
rect 128100 13100 128500 13500
rect 128100 12600 128500 13000
rect 128100 12100 128500 12500
rect 144582 14100 144982 14500
rect 144582 13600 144982 14000
rect 144582 13100 144982 13500
rect 144582 12600 144982 13000
rect 144582 12100 144982 12500
<< metal3 >>
rect 16194 693000 21194 704800
rect 68194 703374 73194 704800
rect 68194 702300 73200 703374
rect 68200 702000 73200 702300
rect 68194 698000 73200 702000
rect 51500 693400 57500 693500
rect 51500 693000 51600 693400
rect 16194 688000 51600 693000
rect 51500 687600 51600 688000
rect 57400 687600 57500 693400
rect 68200 693000 73200 698000
rect 120194 694000 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect 119700 693900 125700 694000
rect 99500 693400 105500 693500
rect 99500 693000 99600 693400
rect 68200 688000 99600 693000
rect 51500 687500 57500 687600
rect 99500 687600 99600 688000
rect 105400 687600 105500 693400
rect 119700 688100 119800 693900
rect 125600 688100 125700 693900
rect 119700 688000 125700 688100
rect 99500 687500 105500 687600
rect 33000 685600 39000 685700
rect 33000 685242 33100 685600
rect -800 680242 33100 685242
rect 33000 679800 33100 680242
rect 38900 685242 39000 685600
rect 38900 680242 39004 685242
rect 38900 679800 39000 680242
rect 33000 679700 39000 679800
rect 582300 677984 584800 682984
rect -800 643842 1660 648642
rect 582340 639784 584800 644584
rect -800 633842 10010 638642
rect 5990 608989 10010 633842
rect 582340 629784 584800 634584
rect 5991 581000 10010 608989
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 16000 582600 24000 583000
rect 16000 581000 16400 582600
rect 5991 577000 16400 581000
rect 5991 576991 10010 577000
rect 16000 575400 16400 577000
rect 23600 575400 24000 582600
rect 16000 575000 24000 575400
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 910 511880 20000 511890
rect 900 511870 20000 511880
rect 890 511860 20000 511870
rect 880 511850 20000 511860
rect 870 511840 20000 511850
rect 860 511830 20000 511840
rect 850 511820 20000 511830
rect 840 511810 20000 511820
rect 830 511800 20000 511810
rect 820 511790 20000 511800
rect 810 511780 20000 511790
rect 800 511770 20000 511780
rect 790 511760 20000 511770
rect 780 511750 20000 511760
rect 770 511740 20000 511750
rect 760 511730 20000 511740
rect 750 511720 20000 511730
rect 740 511710 20000 511720
rect 730 511700 20000 511710
rect 720 511690 20000 511700
rect 710 511680 20000 511690
rect 700 511670 20000 511680
rect 690 511660 20000 511670
rect 680 511650 20000 511660
rect 670 511642 20000 511650
rect -800 511530 20000 511642
rect 670 511520 20000 511530
rect 680 511510 20000 511520
rect 690 511500 20000 511510
rect 700 511490 20000 511500
rect 710 511480 20000 511490
rect 720 511470 20000 511480
rect 730 511460 20000 511470
rect 740 511450 20000 511460
rect 750 511440 20000 511450
rect 760 511430 20000 511440
rect 770 511420 20000 511430
rect 780 511410 20000 511420
rect 790 511400 20000 511410
rect 800 511390 20000 511400
rect 810 511380 20000 511390
rect 820 511370 20000 511380
rect 830 511360 20000 511370
rect 840 511350 20000 511360
rect 850 511340 20000 511350
rect 860 511330 20000 511340
rect 870 511320 20000 511330
rect 880 511310 20000 511320
rect 890 511300 20000 511310
rect 900 511290 20000 511300
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 840 468660 16000 468670
rect 830 468650 16000 468660
rect 820 468640 16000 468650
rect 810 468630 16000 468640
rect 800 468620 16000 468630
rect 790 468610 16000 468620
rect 780 468600 16000 468610
rect 770 468590 16000 468600
rect 760 468580 16000 468590
rect 750 468570 16000 468580
rect 740 468560 16000 468570
rect 730 468550 16000 468560
rect 720 468540 16000 468550
rect 710 468530 16000 468540
rect 700 468520 16000 468530
rect 690 468510 16000 468520
rect 680 468500 16000 468510
rect 670 468490 16000 468500
rect 660 468480 16000 468490
rect 650 468470 16000 468480
rect 640 468460 16000 468470
rect 630 468450 16000 468460
rect 620 468440 16000 468450
rect 610 468430 16000 468440
rect 600 468420 16000 468430
rect -800 468308 16000 468420
rect 600 468300 16000 468308
rect 610 468290 16000 468300
rect 620 468280 16000 468290
rect 630 468270 16000 468280
rect 640 468260 16000 468270
rect 650 468250 16000 468260
rect 660 468240 16000 468250
rect 670 468230 16000 468240
rect 680 468220 16000 468230
rect 690 468210 16000 468220
rect 700 468200 16000 468210
rect 710 468190 16000 468200
rect 720 468180 16000 468190
rect 730 468170 16000 468180
rect 740 468160 16000 468170
rect 750 468150 16000 468160
rect 760 468140 16000 468150
rect 770 468130 16000 468140
rect 780 468120 16000 468130
rect 790 468110 16000 468120
rect 800 468100 16000 468110
rect 810 468090 16000 468100
rect 820 468080 16000 468090
rect 830 468070 16000 468080
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 840 425440 12000 425450
rect 830 425430 12000 425440
rect 820 425420 12000 425430
rect 810 425410 12000 425420
rect 800 425400 12000 425410
rect 790 425390 12000 425400
rect 780 425380 12000 425390
rect 770 425370 12000 425380
rect 760 425360 12000 425370
rect 750 425350 12000 425360
rect 740 425340 12000 425350
rect 730 425330 12000 425340
rect 720 425320 12000 425330
rect 710 425310 12000 425320
rect 700 425300 12000 425310
rect 690 425290 12000 425300
rect 680 425280 12000 425290
rect 670 425270 12000 425280
rect 660 425260 12000 425270
rect 650 425250 12000 425260
rect 640 425240 12000 425250
rect 630 425230 12000 425240
rect 620 425220 12000 425230
rect 610 425210 12000 425220
rect 600 425198 12000 425210
rect -800 425086 12000 425198
rect 600 425080 12000 425086
rect 610 425070 12000 425080
rect 620 425060 12000 425070
rect 630 425050 12000 425060
rect 640 425040 12000 425050
rect 650 425030 12000 425040
rect 660 425020 12000 425030
rect 670 425010 12000 425020
rect 680 425000 12000 425010
rect 690 424990 12000 425000
rect 700 424980 12000 424990
rect 710 424970 12000 424980
rect 720 424960 12000 424970
rect 730 424950 12000 424960
rect 740 424940 12000 424950
rect 750 424930 12000 424940
rect 760 424920 12000 424930
rect 770 424910 12000 424920
rect 780 424900 12000 424910
rect 790 424890 12000 424900
rect 800 424880 12000 424890
rect 810 424870 12000 424880
rect 820 424860 12000 424870
rect 830 424850 12000 424860
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 10000 393160 12000 424850
rect 14000 396795 16000 468070
rect 18000 400284 20000 511290
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 30988 400284 33718 400289
rect 18000 400264 33718 400284
rect 18000 399704 31048 400264
rect 31608 399704 31748 400264
rect 32308 399704 32448 400264
rect 33008 399704 33148 400264
rect 33708 399704 33718 400264
rect 18000 399564 33718 399704
rect 18000 399004 31048 399564
rect 31608 399004 31748 399564
rect 32308 399004 32448 399564
rect 33008 399004 33148 399564
rect 33708 399004 33718 399564
rect 18000 398864 33718 399004
rect 18000 398304 31048 398864
rect 31608 398304 31748 398864
rect 32308 398304 32448 398864
rect 33008 398304 33148 398864
rect 33708 398304 33718 398864
rect 18000 398284 33718 398304
rect 31628 398274 31728 398284
rect 30960 396795 33690 396803
rect 14000 396778 33690 396795
rect 14000 396218 31020 396778
rect 31580 396218 31720 396778
rect 32280 396218 32420 396778
rect 32980 396218 33120 396778
rect 33680 396218 33690 396778
rect 14000 396078 33690 396218
rect 14000 395518 31020 396078
rect 31580 395518 31720 396078
rect 32280 395518 32420 396078
rect 32980 395518 33120 396078
rect 33680 395518 33690 396078
rect 14000 395378 33690 395518
rect 14000 394818 31020 395378
rect 31580 394818 31720 395378
rect 32280 394818 32420 395378
rect 32980 394818 33120 395378
rect 33680 394818 33690 395378
rect 14000 394798 33690 394818
rect 14000 394795 33261 394798
rect 31600 394788 31700 394795
rect 31028 393160 33758 393163
rect 10000 393138 33758 393160
rect 10000 392578 31088 393138
rect 31648 392578 31788 393138
rect 32348 392578 32488 393138
rect 33048 392578 33188 393138
rect 33748 392578 33758 393138
rect 10000 392438 33758 392578
rect 10000 391878 31088 392438
rect 31648 391878 31788 392438
rect 32348 391878 32488 392438
rect 33048 391878 33188 392438
rect 33748 391878 33758 392438
rect 10000 391738 33758 391878
rect 10000 391178 31088 391738
rect 31648 391178 31788 391738
rect 32348 391178 32488 391738
rect 33048 391178 33188 391738
rect 33748 391178 33758 391738
rect 10000 391160 33758 391178
rect 31068 391158 33758 391160
rect 31668 391148 31768 391158
rect 31028 389055 33758 389059
rect 4000 389034 33758 389055
rect 4000 388474 31088 389034
rect 31648 388474 31788 389034
rect 32348 388474 32488 389034
rect 33048 388474 33188 389034
rect 33748 388474 33758 389034
rect 4000 388334 33758 388474
rect 4000 387774 31088 388334
rect 31648 387774 31788 388334
rect 32348 387774 32488 388334
rect 33048 387774 33188 388334
rect 33748 387774 33758 388334
rect 4000 387634 33758 387774
rect 4000 387074 31088 387634
rect 31648 387074 31788 387634
rect 32348 387074 32488 387634
rect 33048 387074 33188 387634
rect 33748 387074 33758 387634
rect 4000 387055 33758 387074
rect 4000 382230 6000 387055
rect 31068 387054 33758 387055
rect 31668 387044 31768 387054
rect 840 382220 6000 382230
rect 830 382210 6000 382220
rect 820 382200 6000 382210
rect 810 382190 6000 382200
rect 800 382180 6000 382190
rect 790 382170 6000 382180
rect 780 382160 6000 382170
rect 770 382150 6000 382160
rect 760 382140 6000 382150
rect 750 382130 6000 382140
rect 740 382120 6000 382130
rect 730 382110 6000 382120
rect 720 382100 6000 382110
rect 710 382090 6000 382100
rect 700 382080 6000 382090
rect 690 382070 6000 382080
rect 680 382060 6000 382070
rect 670 382050 6000 382060
rect 660 382040 6000 382050
rect 650 382030 6000 382040
rect 640 382020 6000 382030
rect 630 382010 6000 382020
rect 620 382000 6000 382010
rect 610 381990 6000 382000
rect 600 381976 6000 381990
rect -800 381864 6000 381976
rect 600 381860 6000 381864
rect 610 381850 6000 381860
rect 620 381840 6000 381850
rect 630 381830 6000 381840
rect 640 381820 6000 381830
rect 650 381810 6000 381820
rect 660 381800 6000 381810
rect 670 381790 6000 381800
rect 680 381780 6000 381790
rect 690 381770 6000 381780
rect 700 381760 6000 381770
rect 710 381750 6000 381760
rect 720 381740 6000 381750
rect 730 381730 6000 381740
rect 740 381720 6000 381730
rect 750 381710 6000 381720
rect 760 381700 6000 381710
rect 770 381690 6000 381700
rect 780 381680 6000 381690
rect 790 381670 6000 381680
rect 800 381660 6000 381670
rect 810 381650 6000 381660
rect 820 381640 6000 381650
rect 830 381630 6000 381640
rect 8000 385590 33890 385615
rect 8000 385030 31220 385590
rect 31780 385030 31920 385590
rect 32480 385030 32620 385590
rect 33180 385030 33320 385590
rect 33880 385030 33890 385590
rect 8000 384890 33890 385030
rect 8000 384330 31220 384890
rect 31780 384330 31920 384890
rect 32480 384330 32620 384890
rect 33180 384330 33320 384890
rect 33880 384330 33890 384890
rect 8000 384190 33890 384330
rect 8000 383630 31220 384190
rect 31780 383630 31920 384190
rect 32480 383630 32620 384190
rect 33180 383630 33320 384190
rect 33880 383630 33890 384190
rect 8000 383615 33890 383630
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 8000 339010 10000 383615
rect 31200 383610 33890 383615
rect 31800 383600 31900 383610
rect 840 339000 10000 339010
rect 830 338990 10000 339000
rect 820 338980 10000 338990
rect 810 338970 10000 338980
rect 800 338960 10000 338970
rect 790 338950 10000 338960
rect 780 338940 10000 338950
rect 770 338930 10000 338940
rect 760 338920 10000 338930
rect 750 338910 10000 338920
rect 740 338900 10000 338910
rect 730 338890 10000 338900
rect 720 338880 10000 338890
rect 710 338870 10000 338880
rect 700 338860 10000 338870
rect 690 338850 10000 338860
rect 680 338840 10000 338850
rect 670 338830 10000 338840
rect 660 338820 10000 338830
rect 650 338810 10000 338820
rect 640 338800 10000 338810
rect 630 338790 10000 338800
rect 620 338780 10000 338790
rect 610 338770 10000 338780
rect 600 338754 10000 338770
rect -800 338642 10000 338754
rect 600 338640 10000 338642
rect 610 338630 10000 338640
rect 620 338620 10000 338630
rect 630 338610 10000 338620
rect 640 338600 10000 338610
rect 650 338590 10000 338600
rect 660 338580 10000 338590
rect 670 338570 10000 338580
rect 680 338560 10000 338570
rect 690 338550 10000 338560
rect 700 338540 10000 338550
rect 710 338530 10000 338540
rect 720 338520 10000 338530
rect 730 338510 10000 338520
rect 740 338500 10000 338510
rect 750 338490 10000 338500
rect 760 338480 10000 338490
rect 770 338470 10000 338480
rect 780 338460 10000 338470
rect 790 338450 10000 338460
rect 800 338440 10000 338450
rect 810 338430 10000 338440
rect 820 338420 10000 338430
rect 830 338410 10000 338420
rect 12000 377571 81364 377580
rect 12000 377271 78504 377571
rect 78804 377271 78864 377571
rect 79164 377271 79224 377571
rect 79524 377271 79584 377571
rect 79884 377271 79944 377571
rect 80244 377271 80304 377571
rect 80604 377271 80664 377571
rect 80964 377271 81024 377571
rect 81324 377271 81364 377571
rect 12000 377211 81364 377271
rect 12000 376911 78504 377211
rect 78804 376911 78864 377211
rect 79164 376911 79224 377211
rect 79524 376911 79584 377211
rect 79884 376911 79944 377211
rect 80244 376911 80304 377211
rect 80604 376911 80664 377211
rect 80964 376911 81024 377211
rect 81324 376911 81364 377211
rect 12000 376851 81364 376911
rect 12000 376551 78504 376851
rect 78804 376551 78864 376851
rect 79164 376551 79224 376851
rect 79524 376551 79584 376851
rect 79884 376551 79944 376851
rect 80244 376551 80304 376851
rect 80604 376551 80664 376851
rect 80964 376551 81024 376851
rect 81324 376551 81364 376851
rect 12000 376491 81364 376551
rect 12000 376191 78504 376491
rect 78804 376191 78864 376491
rect 79164 376191 79224 376491
rect 79524 376191 79584 376491
rect 79884 376191 79944 376491
rect 80244 376191 80304 376491
rect 80604 376191 80664 376491
rect 80964 376191 81024 376491
rect 81324 376191 81364 376491
rect 12000 376131 81364 376191
rect 12000 375831 78504 376131
rect 78804 375831 78864 376131
rect 79164 375831 79224 376131
rect 79524 375831 79584 376131
rect 79884 375831 79944 376131
rect 80244 375831 80304 376131
rect 80604 375831 80664 376131
rect 80964 375831 81024 376131
rect 81324 375831 81364 376131
rect 12000 375771 81364 375831
rect 12000 375580 78504 375771
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 12000 295780 14000 375580
rect 78496 375471 78504 375580
rect 78804 375471 78864 375771
rect 79164 375471 79224 375771
rect 79524 375471 79584 375771
rect 79884 375471 79944 375771
rect 80244 375471 80304 375771
rect 80604 375471 80664 375771
rect 80964 375471 81024 375771
rect 81324 375471 81364 375771
rect 78496 375451 81364 375471
rect 840 295770 14000 295780
rect 830 295760 14000 295770
rect 820 295750 14000 295760
rect 810 295740 14000 295750
rect 800 295730 14000 295740
rect 790 295720 14000 295730
rect 780 295710 14000 295720
rect 770 295700 14000 295710
rect 760 295690 14000 295700
rect 750 295680 14000 295690
rect 740 295670 14000 295680
rect 730 295660 14000 295670
rect 720 295650 14000 295660
rect 710 295640 14000 295650
rect 700 295630 14000 295640
rect 690 295620 14000 295630
rect 680 295610 14000 295620
rect 670 295600 14000 295610
rect 660 295590 14000 295600
rect 650 295580 14000 295590
rect 640 295570 14000 295580
rect 630 295560 14000 295570
rect 620 295550 14000 295560
rect 610 295540 14000 295550
rect 600 295532 14000 295540
rect -800 295420 14000 295532
rect 600 295410 14000 295420
rect 610 295400 14000 295410
rect 620 295390 14000 295400
rect 630 295380 14000 295390
rect 640 295370 14000 295380
rect 650 295360 14000 295370
rect 660 295350 14000 295360
rect 670 295340 14000 295350
rect 680 295330 14000 295340
rect 690 295320 14000 295330
rect 700 295310 14000 295320
rect 710 295300 14000 295310
rect 720 295290 14000 295300
rect 730 295280 14000 295290
rect 740 295270 14000 295280
rect 750 295260 14000 295270
rect 760 295250 14000 295260
rect 770 295240 14000 295250
rect 780 295230 14000 295240
rect 790 295220 14000 295230
rect 800 295210 14000 295220
rect 810 295200 14000 295210
rect 820 295190 14000 295200
rect 830 295180 14000 295190
rect 16000 371880 159760 371889
rect 16000 371580 156900 371880
rect 157200 371580 157260 371880
rect 157560 371580 157620 371880
rect 157920 371580 157980 371880
rect 158280 371580 158340 371880
rect 158640 371580 158700 371880
rect 159000 371580 159060 371880
rect 159360 371580 159420 371880
rect 159720 371580 159760 371880
rect 16000 371520 159760 371580
rect 16000 371220 156900 371520
rect 157200 371220 157260 371520
rect 157560 371220 157620 371520
rect 157920 371220 157980 371520
rect 158280 371220 158340 371520
rect 158640 371220 158700 371520
rect 159000 371220 159060 371520
rect 159360 371220 159420 371520
rect 159720 371220 159760 371520
rect 16000 371160 159760 371220
rect 16000 370860 156900 371160
rect 157200 370860 157260 371160
rect 157560 370860 157620 371160
rect 157920 370860 157980 371160
rect 158280 370860 158340 371160
rect 158640 370860 158700 371160
rect 159000 370860 159060 371160
rect 159360 370860 159420 371160
rect 159720 370860 159760 371160
rect 16000 370800 159760 370860
rect 16000 370500 156900 370800
rect 157200 370500 157260 370800
rect 157560 370500 157620 370800
rect 157920 370500 157980 370800
rect 158280 370500 158340 370800
rect 158640 370500 158700 370800
rect 159000 370500 159060 370800
rect 159360 370500 159420 370800
rect 159720 370500 159760 370800
rect 16000 370440 159760 370500
rect 16000 370140 156900 370440
rect 157200 370140 157260 370440
rect 157560 370140 157620 370440
rect 157920 370140 157980 370440
rect 158280 370140 158340 370440
rect 158640 370140 158700 370440
rect 159000 370140 159060 370440
rect 159360 370140 159420 370440
rect 159720 370140 159760 370440
rect 16000 370080 159760 370140
rect 16000 369889 156900 370080
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 16000 252760 18000 369889
rect 156880 369780 156900 369889
rect 157200 369780 157260 370080
rect 157560 369780 157620 370080
rect 157920 369780 157980 370080
rect 158280 369780 158340 370080
rect 158640 369780 158700 370080
rect 159000 369780 159060 370080
rect 159360 369780 159420 370080
rect 159720 369780 159760 370080
rect 156880 369760 159760 369780
rect 840 252750 18000 252760
rect 830 252740 18000 252750
rect 820 252730 18000 252740
rect 810 252720 18000 252730
rect 800 252710 18000 252720
rect 790 252700 18000 252710
rect 780 252690 18000 252700
rect 770 252680 18000 252690
rect 760 252670 18000 252680
rect 750 252660 18000 252670
rect 740 252650 18000 252660
rect 730 252640 18000 252650
rect 720 252630 18000 252640
rect 710 252620 18000 252630
rect 700 252610 18000 252620
rect 690 252600 18000 252610
rect 680 252590 18000 252600
rect 670 252580 18000 252590
rect 660 252570 18000 252580
rect 650 252560 18000 252570
rect 640 252550 18000 252560
rect 630 252540 18000 252550
rect 620 252530 18000 252540
rect 610 252520 18000 252530
rect 600 252510 18000 252520
rect -800 252398 18000 252510
rect 600 252390 18000 252398
rect 610 252380 18000 252390
rect 620 252370 18000 252380
rect 630 252360 18000 252370
rect 640 252350 18000 252360
rect 650 252340 18000 252350
rect 660 252330 18000 252340
rect 670 252320 18000 252330
rect 680 252310 18000 252320
rect 690 252300 18000 252310
rect 700 252290 18000 252300
rect 710 252280 18000 252290
rect 720 252270 18000 252280
rect 730 252260 18000 252270
rect 740 252250 18000 252260
rect 750 252240 18000 252250
rect 760 252230 18000 252240
rect 770 252220 18000 252230
rect 780 252210 18000 252220
rect 790 252200 18000 252210
rect 800 252190 18000 252200
rect 810 252180 18000 252190
rect 820 252170 18000 252180
rect 830 252160 18000 252170
rect 20000 366414 235582 366423
rect 20000 366114 232722 366414
rect 233022 366114 233082 366414
rect 233382 366114 233442 366414
rect 233742 366114 233802 366414
rect 234102 366114 234162 366414
rect 234462 366114 234522 366414
rect 234822 366114 234882 366414
rect 235182 366114 235242 366414
rect 235542 366114 235582 366414
rect 20000 366054 235582 366114
rect 20000 365754 232722 366054
rect 233022 365754 233082 366054
rect 233382 365754 233442 366054
rect 233742 365754 233802 366054
rect 234102 365754 234162 366054
rect 234462 365754 234522 366054
rect 234822 365754 234882 366054
rect 235182 365754 235242 366054
rect 235542 365754 235582 366054
rect 20000 365694 235582 365754
rect 20000 365394 232722 365694
rect 233022 365394 233082 365694
rect 233382 365394 233442 365694
rect 233742 365394 233802 365694
rect 234102 365394 234162 365694
rect 234462 365394 234522 365694
rect 234822 365394 234882 365694
rect 235182 365394 235242 365694
rect 235542 365394 235582 365694
rect 20000 365334 235582 365394
rect 20000 365034 232722 365334
rect 233022 365034 233082 365334
rect 233382 365034 233442 365334
rect 233742 365034 233802 365334
rect 234102 365034 234162 365334
rect 234462 365034 234522 365334
rect 234822 365034 234882 365334
rect 235182 365034 235242 365334
rect 235542 365034 235582 365334
rect 20000 364974 235582 365034
rect 20000 364674 232722 364974
rect 233022 364674 233082 364974
rect 233382 364674 233442 364974
rect 233742 364674 233802 364974
rect 234102 364674 234162 364974
rect 234462 364674 234522 364974
rect 234822 364674 234882 364974
rect 235182 364674 235242 364974
rect 235542 364674 235582 364974
rect 583520 364784 584800 364896
rect 20000 364614 235582 364674
rect 20000 364423 232722 364614
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect -800 177530 13234 177688
rect -800 177230 8080 177530
rect 8380 177230 8440 177530
rect 8740 177230 8800 177530
rect 9100 177230 9160 177530
rect 9460 177230 9520 177530
rect 9820 177230 9880 177530
rect 10180 177230 10240 177530
rect 10540 177230 10600 177530
rect 10900 177230 10960 177530
rect 11260 177230 11320 177530
rect 11620 177230 11680 177530
rect 11980 177230 13234 177530
rect -800 177170 13234 177230
rect -800 176870 8080 177170
rect 8380 176870 8440 177170
rect 8740 176870 8800 177170
rect 9100 176870 9160 177170
rect 9460 176870 9520 177170
rect 9820 176870 9880 177170
rect 10180 176870 10240 177170
rect 10540 176870 10600 177170
rect 10900 176870 10960 177170
rect 11260 176870 11320 177170
rect 11620 176870 11680 177170
rect 11980 176870 13234 177170
rect -800 176810 13234 176870
rect -800 176510 8080 176810
rect 8380 176510 8440 176810
rect 8740 176510 8800 176810
rect 9100 176510 9160 176810
rect 9460 176510 9520 176810
rect 9820 176510 9880 176810
rect 10180 176510 10240 176810
rect 10540 176510 10600 176810
rect 10900 176510 10960 176810
rect 11260 176510 11320 176810
rect 11620 176510 11680 176810
rect 11980 176510 13234 176810
rect -800 176450 13234 176510
rect -800 176150 8080 176450
rect 8380 176150 8440 176450
rect 8740 176150 8800 176450
rect 9100 176150 9160 176450
rect 9460 176150 9520 176450
rect 9820 176150 9880 176450
rect 10180 176150 10240 176450
rect 10540 176150 10600 176450
rect 10900 176150 10960 176450
rect 11260 176150 11320 176450
rect 11620 176150 11680 176450
rect 11980 176150 13234 176450
rect -800 176090 13234 176150
rect -800 175790 8080 176090
rect 8380 175790 8440 176090
rect 8740 175790 8800 176090
rect 9100 175790 9160 176090
rect 9460 175790 9520 176090
rect 9820 175790 9880 176090
rect 10180 175790 10240 176090
rect 10540 175790 10600 176090
rect 10900 175790 10960 176090
rect 11260 175790 11320 176090
rect 11620 175790 11680 176090
rect 11980 175790 13234 176090
rect -800 175730 13234 175790
rect -800 175430 8080 175730
rect 8380 175430 8440 175730
rect 8740 175430 8800 175730
rect 9100 175430 9160 175730
rect 9460 175430 9520 175730
rect 9820 175430 9880 175730
rect 10180 175430 10240 175730
rect 10540 175430 10600 175730
rect 10900 175430 10960 175730
rect 11260 175430 11320 175730
rect 11620 175430 11680 175730
rect 11980 175430 13234 175730
rect -800 175370 13234 175430
rect -800 175070 8080 175370
rect 8380 175070 8440 175370
rect 8740 175070 8800 175370
rect 9100 175070 9160 175370
rect 9460 175070 9520 175370
rect 9820 175070 9880 175370
rect 10180 175070 10240 175370
rect 10540 175070 10600 175370
rect 10900 175070 10960 175370
rect 11260 175070 11320 175370
rect 11620 175070 11680 175370
rect 11980 175070 13234 175370
rect -800 175010 13234 175070
rect -800 174710 8080 175010
rect 8380 174710 8440 175010
rect 8740 174710 8800 175010
rect 9100 174710 9160 175010
rect 9460 174710 9520 175010
rect 9820 174710 9880 175010
rect 10180 174710 10240 175010
rect 10540 174710 10600 175010
rect 10900 174710 10960 175010
rect 11260 174710 11320 175010
rect 11620 174710 11680 175010
rect 11980 174710 13234 175010
rect -800 174650 13234 174710
rect -800 174350 8080 174650
rect 8380 174350 8440 174650
rect 8740 174350 8800 174650
rect 9100 174350 9160 174650
rect 9460 174350 9520 174650
rect 9820 174350 9880 174650
rect 10180 174350 10240 174650
rect 10540 174350 10600 174650
rect 10900 174350 10960 174650
rect 11260 174350 11320 174650
rect 11620 174350 11680 174650
rect 11980 174350 13234 174650
rect -800 174290 13234 174350
rect -800 173990 8080 174290
rect 8380 173990 8440 174290
rect 8740 173990 8800 174290
rect 9100 173990 9160 174290
rect 9460 173990 9520 174290
rect 9820 173990 9880 174290
rect 10180 173990 10240 174290
rect 10540 173990 10600 174290
rect 10900 173990 10960 174290
rect 11260 173990 11320 174290
rect 11620 173990 11680 174290
rect 11980 173990 13234 174290
rect -800 173930 13234 173990
rect -800 173630 8080 173930
rect 8380 173630 8440 173930
rect 8740 173630 8800 173930
rect 9100 173630 9160 173930
rect 9460 173630 9520 173930
rect 9820 173630 9880 173930
rect 10180 173630 10240 173930
rect 10540 173630 10600 173930
rect 10900 173630 10960 173930
rect 11260 173630 11320 173930
rect 11620 173630 11680 173930
rect 11980 173630 13234 173930
rect -800 173570 13234 173630
rect -800 173270 8080 173570
rect 8380 173270 8440 173570
rect 8740 173270 8800 173570
rect 9100 173270 9160 173570
rect 9460 173270 9520 173570
rect 9820 173270 9880 173570
rect 10180 173270 10240 173570
rect 10540 173270 10600 173570
rect 10900 173270 10960 173570
rect 11260 173270 11320 173570
rect 11620 173270 11680 173570
rect 11980 173270 13234 173570
rect -800 173210 13234 173270
rect -800 172910 8080 173210
rect 8380 172910 8440 173210
rect 8740 172910 8800 173210
rect 9100 172910 9160 173210
rect 9460 172910 9520 173210
rect 9820 172910 9880 173210
rect 10180 172910 10240 173210
rect 10540 172910 10600 173210
rect 10900 172910 10960 173210
rect 11260 172910 11320 173210
rect 11620 172910 11680 173210
rect 11980 172910 13234 173210
rect -800 172888 13234 172910
rect -800 162888 1660 167688
rect 20000 125140 22000 364423
rect 232714 364314 232722 364423
rect 233022 364314 233082 364614
rect 233382 364314 233442 364614
rect 233742 364314 233802 364614
rect 234102 364314 234162 364614
rect 234462 364314 234522 364614
rect 234822 364314 234882 364614
rect 235182 364314 235242 364614
rect 235542 364314 235582 364614
rect 232714 364294 235582 364314
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 840 125130 22000 125140
rect 830 125120 22000 125130
rect 820 125110 22000 125120
rect 810 125100 22000 125110
rect 800 125090 22000 125100
rect 790 125080 22000 125090
rect 780 125070 22000 125080
rect 770 125060 22000 125070
rect 760 125050 22000 125060
rect 750 125040 22000 125050
rect 740 125030 22000 125040
rect 730 125020 22000 125030
rect 720 125010 22000 125020
rect 710 125000 22000 125010
rect 700 124990 22000 125000
rect 690 124980 22000 124990
rect 680 124970 22000 124980
rect 670 124960 22000 124970
rect 660 124950 22000 124960
rect 650 124940 22000 124950
rect 640 124930 22000 124940
rect 630 124920 22000 124930
rect 620 124910 22000 124920
rect 610 124900 22000 124910
rect 600 124888 22000 124900
rect -800 124776 22000 124888
rect 600 124770 22000 124776
rect 610 124760 22000 124770
rect 620 124750 22000 124760
rect 630 124740 22000 124750
rect 640 124730 22000 124740
rect 650 124720 22000 124730
rect 660 124710 22000 124720
rect 670 124700 22000 124710
rect 680 124690 22000 124700
rect 690 124680 22000 124690
rect 700 124670 22000 124680
rect 710 124660 22000 124670
rect 720 124650 22000 124660
rect 730 124640 22000 124650
rect 740 124630 22000 124640
rect 750 124620 22000 124630
rect 760 124610 22000 124620
rect 770 124600 22000 124610
rect 780 124590 22000 124600
rect 790 124580 22000 124590
rect 800 124570 22000 124580
rect 810 124560 22000 124570
rect 820 124550 22000 124560
rect 830 124540 22000 124550
rect 24000 360188 313380 360197
rect 24000 359888 310516 360188
rect 310816 359888 310876 360188
rect 311176 359888 311236 360188
rect 311536 359888 311596 360188
rect 311896 359888 311956 360188
rect 312256 359888 312316 360188
rect 312616 359888 312676 360188
rect 312976 359888 313036 360188
rect 313336 359888 313380 360188
rect 583520 360056 584800 360168
rect 24000 359828 313380 359888
rect 24000 359528 310516 359828
rect 310816 359528 310876 359828
rect 311176 359528 311236 359828
rect 311536 359528 311596 359828
rect 311896 359528 311956 359828
rect 312256 359528 312316 359828
rect 312616 359528 312676 359828
rect 312976 359528 313036 359828
rect 313336 359528 313380 359828
rect 24000 359468 313380 359528
rect 24000 359168 310516 359468
rect 310816 359168 310876 359468
rect 311176 359168 311236 359468
rect 311536 359168 311596 359468
rect 311896 359168 311956 359468
rect 312256 359168 312316 359468
rect 312616 359168 312676 359468
rect 312976 359168 313036 359468
rect 313336 359168 313380 359468
rect 24000 359108 313380 359168
rect 24000 358808 310516 359108
rect 310816 358808 310876 359108
rect 311176 358808 311236 359108
rect 311536 358808 311596 359108
rect 311896 358808 311956 359108
rect 312256 358808 312316 359108
rect 312616 358808 312676 359108
rect 312976 358808 313036 359108
rect 313336 358808 313380 359108
rect 583520 358874 584800 358986
rect 24000 358748 313380 358808
rect 24000 358448 310516 358748
rect 310816 358448 310876 358748
rect 311176 358448 311236 358748
rect 311536 358448 311596 358748
rect 311896 358448 311956 358748
rect 312256 358448 312316 358748
rect 312616 358448 312676 358748
rect 312976 358448 313036 358748
rect 313336 358448 313380 358748
rect 24000 358388 313380 358448
rect 24000 358197 310516 358388
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 24000 81920 26000 358197
rect 310508 358088 310516 358197
rect 310816 358088 310876 358388
rect 311176 358088 311236 358388
rect 311536 358088 311596 358388
rect 311896 358088 311956 358388
rect 312256 358088 312316 358388
rect 312616 358088 312676 358388
rect 312976 358088 313036 358388
rect 313336 358197 313380 358388
rect 313336 358088 313376 358197
rect 310508 358068 313376 358088
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 840 81910 26000 81920
rect 830 81900 26000 81910
rect 820 81890 26000 81900
rect 810 81880 26000 81890
rect 800 81870 26000 81880
rect 790 81860 26000 81870
rect 780 81850 26000 81860
rect 770 81840 26000 81850
rect 760 81830 26000 81840
rect 750 81820 26000 81830
rect 740 81810 26000 81820
rect 730 81800 26000 81810
rect 720 81790 26000 81800
rect 710 81780 26000 81790
rect 700 81770 26000 81780
rect 690 81760 26000 81770
rect 680 81750 26000 81760
rect 670 81740 26000 81750
rect 660 81730 26000 81740
rect 650 81720 26000 81730
rect 640 81710 26000 81720
rect 630 81700 26000 81710
rect 620 81690 26000 81700
rect 610 81680 26000 81690
rect 600 81666 26000 81680
rect -800 81554 26000 81666
rect 600 81550 26000 81554
rect 610 81540 26000 81550
rect 620 81530 26000 81540
rect 630 81520 26000 81530
rect 640 81510 26000 81520
rect 650 81500 26000 81510
rect 660 81490 26000 81500
rect 670 81480 26000 81490
rect 680 81470 26000 81480
rect 690 81460 26000 81470
rect 700 81450 26000 81460
rect 710 81440 26000 81450
rect 720 81430 26000 81440
rect 730 81420 26000 81430
rect 740 81410 26000 81420
rect 750 81400 26000 81410
rect 760 81390 26000 81400
rect 770 81380 26000 81390
rect 780 81370 26000 81380
rect 790 81360 26000 81370
rect 800 81350 26000 81360
rect 810 81340 26000 81350
rect 820 81330 26000 81340
rect 830 81320 26000 81330
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect 840 35140 131200 35150
rect 830 35130 131200 35140
rect 820 35120 131200 35130
rect 810 35110 131200 35120
rect 800 35100 131200 35110
rect 790 35090 131200 35100
rect 780 35080 131200 35090
rect 770 35070 131200 35080
rect 760 35060 131200 35070
rect 750 35050 131200 35060
rect 740 35040 131200 35050
rect 730 35030 131200 35040
rect 720 35020 131200 35030
rect 710 35010 131200 35020
rect 700 35000 131200 35010
rect 690 34990 131200 35000
rect 680 34980 131200 34990
rect 670 34970 131200 34980
rect 660 34960 131200 34970
rect 650 34950 131200 34960
rect 640 34940 131200 34950
rect 630 34930 131200 34940
rect 620 34920 131200 34930
rect 610 34910 131200 34920
rect 600 34898 131200 34910
rect -800 34786 131200 34898
rect 600 34780 131200 34786
rect 610 34770 131200 34780
rect 620 34760 131200 34770
rect 630 34750 131200 34760
rect 640 34740 131200 34750
rect 650 34730 131200 34740
rect 660 34720 131200 34730
rect 670 34710 131200 34720
rect 680 34700 131200 34710
rect 690 34690 131200 34700
rect 700 34680 131200 34690
rect 710 34670 131200 34680
rect 720 34660 131200 34670
rect 730 34650 131200 34660
rect 740 34640 131200 34650
rect 750 34630 131200 34640
rect 760 34620 131200 34630
rect 770 34610 131200 34620
rect 780 34600 131200 34610
rect 790 34590 131200 34600
rect 800 34580 131200 34590
rect 810 34570 131200 34580
rect 820 34560 131200 34570
rect 830 34550 131200 34560
rect 131800 34550 131960 35150
rect 132560 34550 132740 35150
rect 133340 34550 133500 35150
rect 134100 34550 134155 35150
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 110590 15580 110600 16020
rect 111040 15580 111050 16020
rect 114800 15580 114810 16020
rect 115250 15580 115260 16020
rect 119230 15580 119240 16020
rect 119680 15580 119690 16020
rect 123590 15580 123600 16020
rect 124040 15580 124050 16020
rect 128070 15580 128080 16020
rect 128520 15580 128530 16020
rect 583520 15728 584800 15840
rect 110590 15080 110600 15520
rect 111040 15080 111050 15520
rect 114800 15080 114810 15520
rect 115250 15080 115260 15520
rect 119230 15080 119240 15520
rect 119680 15080 119690 15520
rect 123590 15080 123600 15520
rect 124040 15080 124050 15520
rect 128070 15080 128080 15520
rect 128520 15080 128530 15520
rect -800 14546 480 14658
rect 110590 14580 110600 15020
rect 111040 14580 111050 15020
rect 114800 14580 114810 15020
rect 115250 14580 115260 15020
rect 119230 14580 119240 15020
rect 119680 14580 119690 15020
rect 123590 14580 123600 15020
rect 124040 14580 124050 15020
rect 128070 14580 128080 15020
rect 128520 14580 128530 15020
rect 583520 14546 584800 14658
rect 110590 14080 110600 14520
rect 111040 14080 111050 14520
rect 114800 14080 114810 14520
rect 115250 14080 115260 14520
rect 119230 14080 119240 14520
rect 119680 14080 119690 14520
rect 123590 14080 123600 14520
rect 124040 14080 124050 14520
rect 128070 14080 128080 14520
rect 128520 14080 128530 14520
rect 144552 14080 144562 14520
rect 145002 14080 145012 14520
rect 110590 13580 110600 14020
rect 111040 13580 111050 14020
rect 114800 13580 114810 14020
rect 115250 13580 115260 14020
rect 119230 13580 119240 14020
rect 119680 13580 119690 14020
rect 123590 13580 123600 14020
rect 124040 13580 124050 14020
rect 128070 13580 128080 14020
rect 128520 13580 128530 14020
rect 144552 13580 144562 14020
rect 145002 13580 145012 14020
rect -800 13364 480 13476
rect 110590 13080 110600 13520
rect 111040 13080 111050 13520
rect 114800 13080 114810 13520
rect 115250 13080 115260 13520
rect 119230 13080 119240 13520
rect 119680 13080 119690 13520
rect 123590 13080 123600 13520
rect 124040 13080 124050 13520
rect 128070 13080 128080 13520
rect 128520 13080 128530 13520
rect 144552 13080 144562 13520
rect 145002 13080 145012 13520
rect 583520 13364 584800 13476
rect 110590 12580 110600 13020
rect 111040 12580 111050 13020
rect 114800 12580 114810 13020
rect 115250 12580 115260 13020
rect 119230 12580 119240 13020
rect 119680 12580 119690 13020
rect 123590 12580 123600 13020
rect 124040 12580 124050 13020
rect 128070 12580 128080 13020
rect 128520 12580 128530 13020
rect 144552 12580 144562 13020
rect 145002 12580 145012 13020
rect -800 12182 480 12294
rect 110590 12080 110600 12520
rect 111040 12080 111050 12520
rect 114800 12080 114810 12520
rect 115250 12080 115260 12520
rect 119230 12080 119240 12520
rect 119680 12080 119690 12520
rect 123590 12080 123600 12520
rect 124040 12080 124050 12520
rect 128070 12080 128080 12520
rect 128520 12080 128530 12520
rect 144552 12080 144562 12520
rect 145002 12080 145012 12520
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 51600 687600 57400 693400
rect 99600 687600 105400 693400
rect 119800 688100 125600 693900
rect 33100 679800 38900 685600
rect 16400 575400 23600 582600
rect 31048 399704 31608 400264
rect 31748 399704 32308 400264
rect 32448 399704 33008 400264
rect 33148 399704 33708 400264
rect 31048 399004 31608 399564
rect 31748 399004 32308 399564
rect 32448 399004 33008 399564
rect 33148 399004 33708 399564
rect 31048 398304 31608 398864
rect 31748 398304 32308 398864
rect 32448 398304 33008 398864
rect 33148 398304 33708 398864
rect 31020 396218 31580 396778
rect 31720 396218 32280 396778
rect 32420 396218 32980 396778
rect 33120 396218 33680 396778
rect 31020 395518 31580 396078
rect 31720 395518 32280 396078
rect 32420 395518 32980 396078
rect 33120 395518 33680 396078
rect 31020 394818 31580 395378
rect 31720 394818 32280 395378
rect 32420 394818 32980 395378
rect 33120 394818 33680 395378
rect 31088 392578 31648 393138
rect 31788 392578 32348 393138
rect 32488 392578 33048 393138
rect 33188 392578 33748 393138
rect 31088 391878 31648 392438
rect 31788 391878 32348 392438
rect 32488 391878 33048 392438
rect 33188 391878 33748 392438
rect 31088 391178 31648 391738
rect 31788 391178 32348 391738
rect 32488 391178 33048 391738
rect 33188 391178 33748 391738
rect 31088 388474 31648 389034
rect 31788 388474 32348 389034
rect 32488 388474 33048 389034
rect 33188 388474 33748 389034
rect 31088 387774 31648 388334
rect 31788 387774 32348 388334
rect 32488 387774 33048 388334
rect 33188 387774 33748 388334
rect 31088 387074 31648 387634
rect 31788 387074 32348 387634
rect 32488 387074 33048 387634
rect 33188 387074 33748 387634
rect 31220 385030 31780 385590
rect 31920 385030 32480 385590
rect 32620 385030 33180 385590
rect 33320 385030 33880 385590
rect 31220 384330 31780 384890
rect 31920 384330 32480 384890
rect 32620 384330 33180 384890
rect 33320 384330 33880 384890
rect 31220 383630 31780 384190
rect 31920 383630 32480 384190
rect 32620 383630 33180 384190
rect 33320 383630 33880 384190
rect 78504 377271 78804 377571
rect 78864 377271 79164 377571
rect 79224 377271 79524 377571
rect 79584 377271 79884 377571
rect 79944 377271 80244 377571
rect 80304 377271 80604 377571
rect 80664 377271 80964 377571
rect 81024 377271 81324 377571
rect 78504 376911 78804 377211
rect 78864 376911 79164 377211
rect 79224 376911 79524 377211
rect 79584 376911 79884 377211
rect 79944 376911 80244 377211
rect 80304 376911 80604 377211
rect 80664 376911 80964 377211
rect 81024 376911 81324 377211
rect 78504 376551 78804 376851
rect 78864 376551 79164 376851
rect 79224 376551 79524 376851
rect 79584 376551 79884 376851
rect 79944 376551 80244 376851
rect 80304 376551 80604 376851
rect 80664 376551 80964 376851
rect 81024 376551 81324 376851
rect 78504 376191 78804 376491
rect 78864 376191 79164 376491
rect 79224 376191 79524 376491
rect 79584 376191 79884 376491
rect 79944 376191 80244 376491
rect 80304 376191 80604 376491
rect 80664 376191 80964 376491
rect 81024 376191 81324 376491
rect 78504 375831 78804 376131
rect 78864 375831 79164 376131
rect 79224 375831 79524 376131
rect 79584 375831 79884 376131
rect 79944 375831 80244 376131
rect 80304 375831 80604 376131
rect 80664 375831 80964 376131
rect 81024 375831 81324 376131
rect 78504 375471 78804 375771
rect 78864 375471 79164 375771
rect 79224 375471 79524 375771
rect 79584 375471 79884 375771
rect 79944 375471 80244 375771
rect 80304 375471 80604 375771
rect 80664 375471 80964 375771
rect 81024 375471 81324 375771
rect 156900 371580 157200 371880
rect 157260 371580 157560 371880
rect 157620 371580 157920 371880
rect 157980 371580 158280 371880
rect 158340 371580 158640 371880
rect 158700 371580 159000 371880
rect 159060 371580 159360 371880
rect 159420 371580 159720 371880
rect 156900 371220 157200 371520
rect 157260 371220 157560 371520
rect 157620 371220 157920 371520
rect 157980 371220 158280 371520
rect 158340 371220 158640 371520
rect 158700 371220 159000 371520
rect 159060 371220 159360 371520
rect 159420 371220 159720 371520
rect 156900 370860 157200 371160
rect 157260 370860 157560 371160
rect 157620 370860 157920 371160
rect 157980 370860 158280 371160
rect 158340 370860 158640 371160
rect 158700 370860 159000 371160
rect 159060 370860 159360 371160
rect 159420 370860 159720 371160
rect 156900 370500 157200 370800
rect 157260 370500 157560 370800
rect 157620 370500 157920 370800
rect 157980 370500 158280 370800
rect 158340 370500 158640 370800
rect 158700 370500 159000 370800
rect 159060 370500 159360 370800
rect 159420 370500 159720 370800
rect 156900 370140 157200 370440
rect 157260 370140 157560 370440
rect 157620 370140 157920 370440
rect 157980 370140 158280 370440
rect 158340 370140 158640 370440
rect 158700 370140 159000 370440
rect 159060 370140 159360 370440
rect 159420 370140 159720 370440
rect 156900 369780 157200 370080
rect 157260 369780 157560 370080
rect 157620 369780 157920 370080
rect 157980 369780 158280 370080
rect 158340 369780 158640 370080
rect 158700 369780 159000 370080
rect 159060 369780 159360 370080
rect 159420 369780 159720 370080
rect 232722 366114 233022 366414
rect 233082 366114 233382 366414
rect 233442 366114 233742 366414
rect 233802 366114 234102 366414
rect 234162 366114 234462 366414
rect 234522 366114 234822 366414
rect 234882 366114 235182 366414
rect 235242 366114 235542 366414
rect 232722 365754 233022 366054
rect 233082 365754 233382 366054
rect 233442 365754 233742 366054
rect 233802 365754 234102 366054
rect 234162 365754 234462 366054
rect 234522 365754 234822 366054
rect 234882 365754 235182 366054
rect 235242 365754 235542 366054
rect 232722 365394 233022 365694
rect 233082 365394 233382 365694
rect 233442 365394 233742 365694
rect 233802 365394 234102 365694
rect 234162 365394 234462 365694
rect 234522 365394 234822 365694
rect 234882 365394 235182 365694
rect 235242 365394 235542 365694
rect 232722 365034 233022 365334
rect 233082 365034 233382 365334
rect 233442 365034 233742 365334
rect 233802 365034 234102 365334
rect 234162 365034 234462 365334
rect 234522 365034 234822 365334
rect 234882 365034 235182 365334
rect 235242 365034 235542 365334
rect 232722 364674 233022 364974
rect 233082 364674 233382 364974
rect 233442 364674 233742 364974
rect 233802 364674 234102 364974
rect 234162 364674 234462 364974
rect 234522 364674 234822 364974
rect 234882 364674 235182 364974
rect 235242 364674 235542 364974
rect 8080 177230 8380 177530
rect 8440 177230 8740 177530
rect 8800 177230 9100 177530
rect 9160 177230 9460 177530
rect 9520 177230 9820 177530
rect 9880 177230 10180 177530
rect 10240 177230 10540 177530
rect 10600 177230 10900 177530
rect 10960 177230 11260 177530
rect 11320 177230 11620 177530
rect 11680 177230 11980 177530
rect 8080 176870 8380 177170
rect 8440 176870 8740 177170
rect 8800 176870 9100 177170
rect 9160 176870 9460 177170
rect 9520 176870 9820 177170
rect 9880 176870 10180 177170
rect 10240 176870 10540 177170
rect 10600 176870 10900 177170
rect 10960 176870 11260 177170
rect 11320 176870 11620 177170
rect 11680 176870 11980 177170
rect 8080 176510 8380 176810
rect 8440 176510 8740 176810
rect 8800 176510 9100 176810
rect 9160 176510 9460 176810
rect 9520 176510 9820 176810
rect 9880 176510 10180 176810
rect 10240 176510 10540 176810
rect 10600 176510 10900 176810
rect 10960 176510 11260 176810
rect 11320 176510 11620 176810
rect 11680 176510 11980 176810
rect 8080 176150 8380 176450
rect 8440 176150 8740 176450
rect 8800 176150 9100 176450
rect 9160 176150 9460 176450
rect 9520 176150 9820 176450
rect 9880 176150 10180 176450
rect 10240 176150 10540 176450
rect 10600 176150 10900 176450
rect 10960 176150 11260 176450
rect 11320 176150 11620 176450
rect 11680 176150 11980 176450
rect 8080 175790 8380 176090
rect 8440 175790 8740 176090
rect 8800 175790 9100 176090
rect 9160 175790 9460 176090
rect 9520 175790 9820 176090
rect 9880 175790 10180 176090
rect 10240 175790 10540 176090
rect 10600 175790 10900 176090
rect 10960 175790 11260 176090
rect 11320 175790 11620 176090
rect 11680 175790 11980 176090
rect 8080 175430 8380 175730
rect 8440 175430 8740 175730
rect 8800 175430 9100 175730
rect 9160 175430 9460 175730
rect 9520 175430 9820 175730
rect 9880 175430 10180 175730
rect 10240 175430 10540 175730
rect 10600 175430 10900 175730
rect 10960 175430 11260 175730
rect 11320 175430 11620 175730
rect 11680 175430 11980 175730
rect 8080 175070 8380 175370
rect 8440 175070 8740 175370
rect 8800 175070 9100 175370
rect 9160 175070 9460 175370
rect 9520 175070 9820 175370
rect 9880 175070 10180 175370
rect 10240 175070 10540 175370
rect 10600 175070 10900 175370
rect 10960 175070 11260 175370
rect 11320 175070 11620 175370
rect 11680 175070 11980 175370
rect 8080 174710 8380 175010
rect 8440 174710 8740 175010
rect 8800 174710 9100 175010
rect 9160 174710 9460 175010
rect 9520 174710 9820 175010
rect 9880 174710 10180 175010
rect 10240 174710 10540 175010
rect 10600 174710 10900 175010
rect 10960 174710 11260 175010
rect 11320 174710 11620 175010
rect 11680 174710 11980 175010
rect 8080 174350 8380 174650
rect 8440 174350 8740 174650
rect 8800 174350 9100 174650
rect 9160 174350 9460 174650
rect 9520 174350 9820 174650
rect 9880 174350 10180 174650
rect 10240 174350 10540 174650
rect 10600 174350 10900 174650
rect 10960 174350 11260 174650
rect 11320 174350 11620 174650
rect 11680 174350 11980 174650
rect 8080 173990 8380 174290
rect 8440 173990 8740 174290
rect 8800 173990 9100 174290
rect 9160 173990 9460 174290
rect 9520 173990 9820 174290
rect 9880 173990 10180 174290
rect 10240 173990 10540 174290
rect 10600 173990 10900 174290
rect 10960 173990 11260 174290
rect 11320 173990 11620 174290
rect 11680 173990 11980 174290
rect 8080 173630 8380 173930
rect 8440 173630 8740 173930
rect 8800 173630 9100 173930
rect 9160 173630 9460 173930
rect 9520 173630 9820 173930
rect 9880 173630 10180 173930
rect 10240 173630 10540 173930
rect 10600 173630 10900 173930
rect 10960 173630 11260 173930
rect 11320 173630 11620 173930
rect 11680 173630 11980 173930
rect 8080 173270 8380 173570
rect 8440 173270 8740 173570
rect 8800 173270 9100 173570
rect 9160 173270 9460 173570
rect 9520 173270 9820 173570
rect 9880 173270 10180 173570
rect 10240 173270 10540 173570
rect 10600 173270 10900 173570
rect 10960 173270 11260 173570
rect 11320 173270 11620 173570
rect 11680 173270 11980 173570
rect 8080 172910 8380 173210
rect 8440 172910 8740 173210
rect 8800 172910 9100 173210
rect 9160 172910 9460 173210
rect 9520 172910 9820 173210
rect 9880 172910 10180 173210
rect 10240 172910 10540 173210
rect 10600 172910 10900 173210
rect 10960 172910 11260 173210
rect 11320 172910 11620 173210
rect 11680 172910 11980 173210
rect 232722 364314 233022 364614
rect 233082 364314 233382 364614
rect 233442 364314 233742 364614
rect 233802 364314 234102 364614
rect 234162 364314 234462 364614
rect 234522 364314 234822 364614
rect 234882 364314 235182 364614
rect 235242 364314 235542 364614
rect 310516 359888 310816 360188
rect 310876 359888 311176 360188
rect 311236 359888 311536 360188
rect 311596 359888 311896 360188
rect 311956 359888 312256 360188
rect 312316 359888 312616 360188
rect 312676 359888 312976 360188
rect 313036 359888 313336 360188
rect 310516 359528 310816 359828
rect 310876 359528 311176 359828
rect 311236 359528 311536 359828
rect 311596 359528 311896 359828
rect 311956 359528 312256 359828
rect 312316 359528 312616 359828
rect 312676 359528 312976 359828
rect 313036 359528 313336 359828
rect 310516 359168 310816 359468
rect 310876 359168 311176 359468
rect 311236 359168 311536 359468
rect 311596 359168 311896 359468
rect 311956 359168 312256 359468
rect 312316 359168 312616 359468
rect 312676 359168 312976 359468
rect 313036 359168 313336 359468
rect 310516 358808 310816 359108
rect 310876 358808 311176 359108
rect 311236 358808 311536 359108
rect 311596 358808 311896 359108
rect 311956 358808 312256 359108
rect 312316 358808 312616 359108
rect 312676 358808 312976 359108
rect 313036 358808 313336 359108
rect 310516 358448 310816 358748
rect 310876 358448 311176 358748
rect 311236 358448 311536 358748
rect 311596 358448 311896 358748
rect 311956 358448 312256 358748
rect 312316 358448 312616 358748
rect 312676 358448 312976 358748
rect 313036 358448 313336 358748
rect 310516 358088 310816 358388
rect 310876 358088 311176 358388
rect 311236 358088 311536 358388
rect 311596 358088 311896 358388
rect 311956 358088 312256 358388
rect 312316 358088 312616 358388
rect 312676 358088 312976 358388
rect 313036 358088 313336 358388
rect 131200 34550 131800 35150
rect 131960 34550 132560 35150
rect 132740 34550 133340 35150
rect 133500 34550 134100 35150
rect 110600 16000 111040 16020
rect 110600 15600 110620 16000
rect 110620 15600 111020 16000
rect 111020 15600 111040 16000
rect 110600 15580 111040 15600
rect 114810 16000 115250 16020
rect 114810 15600 114830 16000
rect 114830 15600 115230 16000
rect 115230 15600 115250 16000
rect 114810 15580 115250 15600
rect 119240 16000 119680 16020
rect 119240 15600 119260 16000
rect 119260 15600 119660 16000
rect 119660 15600 119680 16000
rect 119240 15580 119680 15600
rect 123600 16000 124040 16020
rect 123600 15600 123620 16000
rect 123620 15600 124020 16000
rect 124020 15600 124040 16000
rect 123600 15580 124040 15600
rect 128080 16000 128520 16020
rect 128080 15600 128100 16000
rect 128100 15600 128500 16000
rect 128500 15600 128520 16000
rect 128080 15580 128520 15600
rect 110600 15500 111040 15520
rect 110600 15100 110620 15500
rect 110620 15100 111020 15500
rect 111020 15100 111040 15500
rect 110600 15080 111040 15100
rect 114810 15500 115250 15520
rect 114810 15100 114830 15500
rect 114830 15100 115230 15500
rect 115230 15100 115250 15500
rect 114810 15080 115250 15100
rect 119240 15500 119680 15520
rect 119240 15100 119260 15500
rect 119260 15100 119660 15500
rect 119660 15100 119680 15500
rect 119240 15080 119680 15100
rect 123600 15500 124040 15520
rect 123600 15100 123620 15500
rect 123620 15100 124020 15500
rect 124020 15100 124040 15500
rect 123600 15080 124040 15100
rect 128080 15500 128520 15520
rect 128080 15100 128100 15500
rect 128100 15100 128500 15500
rect 128500 15100 128520 15500
rect 128080 15080 128520 15100
rect 110600 15000 111040 15020
rect 110600 14600 110620 15000
rect 110620 14600 111020 15000
rect 111020 14600 111040 15000
rect 110600 14580 111040 14600
rect 114810 15000 115250 15020
rect 114810 14600 114830 15000
rect 114830 14600 115230 15000
rect 115230 14600 115250 15000
rect 114810 14580 115250 14600
rect 119240 15000 119680 15020
rect 119240 14600 119260 15000
rect 119260 14600 119660 15000
rect 119660 14600 119680 15000
rect 119240 14580 119680 14600
rect 123600 15000 124040 15020
rect 123600 14600 123620 15000
rect 123620 14600 124020 15000
rect 124020 14600 124040 15000
rect 123600 14580 124040 14600
rect 128080 15000 128520 15020
rect 128080 14600 128100 15000
rect 128100 14600 128500 15000
rect 128500 14600 128520 15000
rect 128080 14580 128520 14600
rect 110600 14500 111040 14520
rect 110600 14100 110620 14500
rect 110620 14100 111020 14500
rect 111020 14100 111040 14500
rect 110600 14080 111040 14100
rect 114810 14500 115250 14520
rect 114810 14100 114830 14500
rect 114830 14100 115230 14500
rect 115230 14100 115250 14500
rect 114810 14080 115250 14100
rect 119240 14500 119680 14520
rect 119240 14100 119260 14500
rect 119260 14100 119660 14500
rect 119660 14100 119680 14500
rect 119240 14080 119680 14100
rect 123600 14500 124040 14520
rect 123600 14100 123620 14500
rect 123620 14100 124020 14500
rect 124020 14100 124040 14500
rect 123600 14080 124040 14100
rect 128080 14500 128520 14520
rect 128080 14100 128100 14500
rect 128100 14100 128500 14500
rect 128500 14100 128520 14500
rect 128080 14080 128520 14100
rect 144562 14500 145002 14520
rect 144562 14100 144582 14500
rect 144582 14100 144982 14500
rect 144982 14100 145002 14500
rect 144562 14080 145002 14100
rect 110600 14000 111040 14020
rect 110600 13600 110620 14000
rect 110620 13600 111020 14000
rect 111020 13600 111040 14000
rect 110600 13580 111040 13600
rect 114810 14000 115250 14020
rect 114810 13600 114830 14000
rect 114830 13600 115230 14000
rect 115230 13600 115250 14000
rect 114810 13580 115250 13600
rect 119240 14000 119680 14020
rect 119240 13600 119260 14000
rect 119260 13600 119660 14000
rect 119660 13600 119680 14000
rect 119240 13580 119680 13600
rect 123600 14000 124040 14020
rect 123600 13600 123620 14000
rect 123620 13600 124020 14000
rect 124020 13600 124040 14000
rect 123600 13580 124040 13600
rect 128080 14000 128520 14020
rect 128080 13600 128100 14000
rect 128100 13600 128500 14000
rect 128500 13600 128520 14000
rect 128080 13580 128520 13600
rect 144562 14000 145002 14020
rect 144562 13600 144582 14000
rect 144582 13600 144982 14000
rect 144982 13600 145002 14000
rect 144562 13580 145002 13600
rect 110600 13500 111040 13520
rect 110600 13100 110620 13500
rect 110620 13100 111020 13500
rect 111020 13100 111040 13500
rect 110600 13080 111040 13100
rect 114810 13500 115250 13520
rect 114810 13100 114830 13500
rect 114830 13100 115230 13500
rect 115230 13100 115250 13500
rect 114810 13080 115250 13100
rect 119240 13500 119680 13520
rect 119240 13100 119260 13500
rect 119260 13100 119660 13500
rect 119660 13100 119680 13500
rect 119240 13080 119680 13100
rect 123600 13500 124040 13520
rect 123600 13100 123620 13500
rect 123620 13100 124020 13500
rect 124020 13100 124040 13500
rect 123600 13080 124040 13100
rect 128080 13500 128520 13520
rect 128080 13100 128100 13500
rect 128100 13100 128500 13500
rect 128500 13100 128520 13500
rect 128080 13080 128520 13100
rect 144562 13500 145002 13520
rect 144562 13100 144582 13500
rect 144582 13100 144982 13500
rect 144982 13100 145002 13500
rect 144562 13080 145002 13100
rect 110600 13000 111040 13020
rect 110600 12600 110620 13000
rect 110620 12600 111020 13000
rect 111020 12600 111040 13000
rect 110600 12580 111040 12600
rect 114810 13000 115250 13020
rect 114810 12600 114830 13000
rect 114830 12600 115230 13000
rect 115230 12600 115250 13000
rect 114810 12580 115250 12600
rect 119240 13000 119680 13020
rect 119240 12600 119260 13000
rect 119260 12600 119660 13000
rect 119660 12600 119680 13000
rect 119240 12580 119680 12600
rect 123600 13000 124040 13020
rect 123600 12600 123620 13000
rect 123620 12600 124020 13000
rect 124020 12600 124040 13000
rect 123600 12580 124040 12600
rect 128080 13000 128520 13020
rect 128080 12600 128100 13000
rect 128100 12600 128500 13000
rect 128500 12600 128520 13000
rect 128080 12580 128520 12600
rect 144562 13000 145002 13020
rect 144562 12600 144582 13000
rect 144582 12600 144982 13000
rect 144982 12600 145002 13000
rect 144562 12580 145002 12600
rect 110600 12500 111040 12520
rect 110600 12100 110620 12500
rect 110620 12100 111020 12500
rect 111020 12100 111040 12500
rect 110600 12080 111040 12100
rect 114810 12500 115250 12520
rect 114810 12100 114830 12500
rect 114830 12100 115230 12500
rect 115230 12100 115250 12500
rect 114810 12080 115250 12100
rect 119240 12500 119680 12520
rect 119240 12100 119260 12500
rect 119260 12100 119660 12500
rect 119660 12100 119680 12500
rect 119240 12080 119680 12100
rect 123600 12500 124040 12520
rect 123600 12100 123620 12500
rect 123620 12100 124020 12500
rect 124020 12100 124040 12500
rect 123600 12080 124040 12100
rect 128080 12500 128520 12520
rect 128080 12100 128100 12500
rect 128100 12100 128500 12500
rect 128500 12100 128520 12500
rect 128080 12080 128520 12100
rect 144562 12500 145002 12520
rect 144562 12100 144582 12500
rect 144582 12100 144982 12500
rect 144982 12100 145002 12500
rect 144562 12080 145002 12100
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 119700 693900 125700 694000
rect 51500 693400 57500 693500
rect 51500 687600 51600 693400
rect 57400 687600 57500 693400
rect 51500 687500 57500 687600
rect 99500 693400 105500 693500
rect 99500 687600 99600 693400
rect 105400 687600 105500 693400
rect 119700 688100 119800 693900
rect 125600 688100 125700 693900
rect 119700 688000 125700 688100
rect 99500 687500 105500 687600
rect 33000 685600 39000 685700
rect 33000 679800 33100 685600
rect 38900 679800 39000 685600
rect 33000 679700 39000 679800
rect 34000 594000 38000 679700
rect 52000 597000 57000 687500
rect 100000 609000 105000 687500
rect 120194 621000 125194 688000
rect 120194 616000 270500 621000
rect 100000 604000 192500 609000
rect 34490 586357 37368 594000
rect 52000 592000 116000 597000
rect 187500 593500 192500 604000
rect 265508 593508 270493 616000
rect 112950 586709 115828 592000
rect 188770 587473 191648 593500
rect 266504 588412 269382 593508
rect 16000 582800 24000 583000
rect 16000 575200 16200 582800
rect 23800 575200 24000 582800
rect 16000 575000 24000 575200
rect 16000 565800 24000 566000
rect 16000 564000 16200 565800
rect 8000 560000 16200 564000
rect 8000 177530 12000 560000
rect 16000 558200 16200 560000
rect 23800 558200 24000 565800
rect 16000 558000 24000 558200
rect 109388 424940 112268 425000
rect 109388 424640 109480 424940
rect 109780 424640 109880 424940
rect 110180 424640 110280 424940
rect 110580 424640 110680 424940
rect 110980 424640 111080 424940
rect 111380 424640 111480 424940
rect 111780 424640 111880 424940
rect 112180 424640 112268 424940
rect 109388 424540 112268 424640
rect 109388 424240 109480 424540
rect 109780 424240 109880 424540
rect 110180 424240 110280 424540
rect 110580 424240 110680 424540
rect 110980 424240 111080 424540
rect 111380 424240 111480 424540
rect 111780 424240 111880 424540
rect 112180 424240 112268 424540
rect 109388 424140 112268 424240
rect 109388 423840 109480 424140
rect 109780 423840 109880 424140
rect 110180 423840 110280 424140
rect 110580 423840 110680 424140
rect 110980 423840 111080 424140
rect 111380 423840 111480 424140
rect 111780 423840 111880 424140
rect 112180 423840 112268 424140
rect 109388 423740 112268 423840
rect 109388 423440 109480 423740
rect 109780 423440 109880 423740
rect 110180 423440 110280 423740
rect 110580 423440 110680 423740
rect 110980 423440 111080 423740
rect 111380 423440 111480 423740
rect 111780 423440 111880 423740
rect 112180 423440 112268 423740
rect 109388 423340 112268 423440
rect 109388 423040 109480 423340
rect 109780 423040 109880 423340
rect 110180 423040 110280 423340
rect 110580 423040 110680 423340
rect 110980 423040 111080 423340
rect 111380 423040 111480 423340
rect 111780 423040 111880 423340
rect 112180 423040 112268 423340
rect 30988 400274 33768 400314
rect 30988 399674 31028 400274
rect 31628 399674 31728 400274
rect 32328 399674 32428 400274
rect 33028 399674 33128 400274
rect 33728 399674 33768 400274
rect 30988 399574 33768 399674
rect 30988 398974 31028 399574
rect 31628 398974 31728 399574
rect 32328 398974 32428 399574
rect 33028 398974 33128 399574
rect 33728 398974 33768 399574
rect 30988 398874 33768 398974
rect 30988 398274 31028 398874
rect 31628 398274 31728 398874
rect 32328 398274 32428 398874
rect 33028 398274 33128 398874
rect 33728 398274 33768 398874
rect 30988 398244 33768 398274
rect 30960 396788 33740 396828
rect 30960 396188 31000 396788
rect 31600 396188 31700 396788
rect 32300 396188 32400 396788
rect 33000 396188 33100 396788
rect 33700 396188 33740 396788
rect 30960 396088 33740 396188
rect 30960 395488 31000 396088
rect 31600 395488 31700 396088
rect 32300 395488 32400 396088
rect 33000 395488 33100 396088
rect 33700 395488 33740 396088
rect 30960 395388 33740 395488
rect 30960 394788 31000 395388
rect 31600 394788 31700 395388
rect 32300 394788 32400 395388
rect 33000 394788 33100 395388
rect 33700 394788 33740 395388
rect 30960 394758 33740 394788
rect 31028 393148 33808 393188
rect 31028 392548 31068 393148
rect 31668 392548 31768 393148
rect 32368 392548 32468 393148
rect 33068 392548 33168 393148
rect 33768 392548 33808 393148
rect 31028 392448 33808 392548
rect 31028 391848 31068 392448
rect 31668 391848 31768 392448
rect 32368 391848 32468 392448
rect 33068 391848 33168 392448
rect 33768 391848 33808 392448
rect 31028 391748 33808 391848
rect 31028 391148 31068 391748
rect 31668 391148 31768 391748
rect 32368 391148 32468 391748
rect 33068 391148 33168 391748
rect 33768 391148 33808 391748
rect 31028 391118 33808 391148
rect 31028 389044 33808 389084
rect 31028 388444 31068 389044
rect 31668 388444 31768 389044
rect 32368 388444 32468 389044
rect 33068 388444 33168 389044
rect 33768 388444 33808 389044
rect 31028 388344 33808 388444
rect 31028 387744 31068 388344
rect 31668 387744 31768 388344
rect 32368 387744 32468 388344
rect 33068 387744 33168 388344
rect 33768 387744 33808 388344
rect 31028 387644 33808 387744
rect 31028 387044 31068 387644
rect 31668 387044 31768 387644
rect 32368 387044 32468 387644
rect 33068 387044 33168 387644
rect 33768 387044 33808 387644
rect 31028 387014 33808 387044
rect 31160 385600 33940 385640
rect 31160 385000 31200 385600
rect 31800 385000 31900 385600
rect 32500 385000 32600 385600
rect 33200 385000 33300 385600
rect 33900 385000 33940 385600
rect 31160 384900 33940 385000
rect 31160 384300 31200 384900
rect 31800 384300 31900 384900
rect 32500 384300 32600 384900
rect 33200 384300 33300 384900
rect 33900 384300 33940 384900
rect 31160 384200 33940 384300
rect 31160 383600 31200 384200
rect 31800 383600 31900 384200
rect 32500 383600 32600 384200
rect 33200 383600 33300 384200
rect 33900 383600 33940 384200
rect 31160 383570 33940 383600
rect 78496 377571 81354 383874
rect 78496 377271 78504 377571
rect 78804 377271 78864 377571
rect 79164 377271 79224 377571
rect 79524 377271 79584 377571
rect 79884 377271 79944 377571
rect 80244 377271 80304 377571
rect 80604 377271 80664 377571
rect 80964 377271 81024 377571
rect 81324 377271 81354 377571
rect 78496 377211 81354 377271
rect 78496 376911 78504 377211
rect 78804 376911 78864 377211
rect 79164 376911 79224 377211
rect 79524 376911 79584 377211
rect 79884 376911 79944 377211
rect 80244 376911 80304 377211
rect 80604 376911 80664 377211
rect 80964 376911 81024 377211
rect 81324 376911 81354 377211
rect 78496 376851 81354 376911
rect 78496 376551 78504 376851
rect 78804 376551 78864 376851
rect 79164 376551 79224 376851
rect 79524 376551 79584 376851
rect 79884 376551 79944 376851
rect 80244 376551 80304 376851
rect 80604 376551 80664 376851
rect 80964 376551 81024 376851
rect 81324 376551 81354 376851
rect 78496 376491 81354 376551
rect 78496 376191 78504 376491
rect 78804 376191 78864 376491
rect 79164 376191 79224 376491
rect 79524 376191 79584 376491
rect 79884 376191 79944 376491
rect 80244 376191 80304 376491
rect 80604 376191 80664 376491
rect 80964 376191 81024 376491
rect 81324 376191 81354 376491
rect 78496 376131 81354 376191
rect 78496 375831 78504 376131
rect 78804 375831 78864 376131
rect 79164 375831 79224 376131
rect 79524 375831 79584 376131
rect 79884 375831 79944 376131
rect 80244 375831 80304 376131
rect 80604 375831 80664 376131
rect 80964 375831 81024 376131
rect 81324 375831 81354 376131
rect 78496 375771 81354 375831
rect 78496 375471 78504 375771
rect 78804 375471 78864 375771
rect 79164 375471 79224 375771
rect 79524 375471 79584 375771
rect 79884 375471 79944 375771
rect 80244 375471 80304 375771
rect 80604 375471 80664 375771
rect 80964 375471 81024 375771
rect 81324 375471 81354 375771
rect 78496 375440 81354 375471
rect 8000 177230 8080 177530
rect 8380 177230 8440 177530
rect 8740 177230 8800 177530
rect 9100 177230 9160 177530
rect 9460 177230 9520 177530
rect 9820 177230 9880 177530
rect 10180 177230 10240 177530
rect 10540 177230 10600 177530
rect 10900 177230 10960 177530
rect 11260 177230 11320 177530
rect 11620 177230 11680 177530
rect 11980 177230 12000 177530
rect 8000 177170 12000 177230
rect 8000 176870 8080 177170
rect 8380 176870 8440 177170
rect 8740 176870 8800 177170
rect 9100 176870 9160 177170
rect 9460 176870 9520 177170
rect 9820 176870 9880 177170
rect 10180 176870 10240 177170
rect 10540 176870 10600 177170
rect 10900 176870 10960 177170
rect 11260 176870 11320 177170
rect 11620 176870 11680 177170
rect 11980 176870 12000 177170
rect 8000 176810 12000 176870
rect 8000 176510 8080 176810
rect 8380 176510 8440 176810
rect 8740 176510 8800 176810
rect 9100 176510 9160 176810
rect 9460 176510 9520 176810
rect 9820 176510 9880 176810
rect 10180 176510 10240 176810
rect 10540 176510 10600 176810
rect 10900 176510 10960 176810
rect 11260 176510 11320 176810
rect 11620 176510 11680 176810
rect 11980 176510 12000 176810
rect 8000 176450 12000 176510
rect 8000 176150 8080 176450
rect 8380 176150 8440 176450
rect 8740 176150 8800 176450
rect 9100 176150 9160 176450
rect 9460 176150 9520 176450
rect 9820 176150 9880 176450
rect 10180 176150 10240 176450
rect 10540 176150 10600 176450
rect 10900 176150 10960 176450
rect 11260 176150 11320 176450
rect 11620 176150 11680 176450
rect 11980 176150 12000 176450
rect 8000 176090 12000 176150
rect 8000 175790 8080 176090
rect 8380 175790 8440 176090
rect 8740 175790 8800 176090
rect 9100 175790 9160 176090
rect 9460 175790 9520 176090
rect 9820 175790 9880 176090
rect 10180 175790 10240 176090
rect 10540 175790 10600 176090
rect 10900 175790 10960 176090
rect 11260 175790 11320 176090
rect 11620 175790 11680 176090
rect 11980 175790 12000 176090
rect 8000 175730 12000 175790
rect 8000 175430 8080 175730
rect 8380 175430 8440 175730
rect 8740 175430 8800 175730
rect 9100 175430 9160 175730
rect 9460 175430 9520 175730
rect 9820 175430 9880 175730
rect 10180 175430 10240 175730
rect 10540 175430 10600 175730
rect 10900 175430 10960 175730
rect 11260 175430 11320 175730
rect 11620 175430 11680 175730
rect 11980 175430 12000 175730
rect 8000 175370 12000 175430
rect 8000 175070 8080 175370
rect 8380 175070 8440 175370
rect 8740 175070 8800 175370
rect 9100 175070 9160 175370
rect 9460 175070 9520 175370
rect 9820 175070 9880 175370
rect 10180 175070 10240 175370
rect 10540 175070 10600 175370
rect 10900 175070 10960 175370
rect 11260 175070 11320 175370
rect 11620 175070 11680 175370
rect 11980 175070 12000 175370
rect 8000 175010 12000 175070
rect 8000 174710 8080 175010
rect 8380 174710 8440 175010
rect 8740 174710 8800 175010
rect 9100 174710 9160 175010
rect 9460 174710 9520 175010
rect 9820 174710 9880 175010
rect 10180 174710 10240 175010
rect 10540 174710 10600 175010
rect 10900 174710 10960 175010
rect 11260 174710 11320 175010
rect 11620 174710 11680 175010
rect 11980 174710 12000 175010
rect 8000 174650 12000 174710
rect 8000 174350 8080 174650
rect 8380 174350 8440 174650
rect 8740 174350 8800 174650
rect 9100 174350 9160 174650
rect 9460 174350 9520 174650
rect 9820 174350 9880 174650
rect 10180 174350 10240 174650
rect 10540 174350 10600 174650
rect 10900 174350 10960 174650
rect 11260 174350 11320 174650
rect 11620 174350 11680 174650
rect 11980 174350 12000 174650
rect 8000 174290 12000 174350
rect 8000 173990 8080 174290
rect 8380 173990 8440 174290
rect 8740 173990 8800 174290
rect 9100 173990 9160 174290
rect 9460 173990 9520 174290
rect 9820 173990 9880 174290
rect 10180 173990 10240 174290
rect 10540 173990 10600 174290
rect 10900 173990 10960 174290
rect 11260 173990 11320 174290
rect 11620 173990 11680 174290
rect 11980 173990 12000 174290
rect 8000 173930 12000 173990
rect 8000 173630 8080 173930
rect 8380 173630 8440 173930
rect 8740 173630 8800 173930
rect 9100 173630 9160 173930
rect 9460 173630 9520 173930
rect 9820 173630 9880 173930
rect 10180 173630 10240 173930
rect 10540 173630 10600 173930
rect 10900 173630 10960 173930
rect 11260 173630 11320 173930
rect 11620 173630 11680 173930
rect 11980 173630 12000 173930
rect 8000 173570 12000 173630
rect 8000 173270 8080 173570
rect 8380 173270 8440 173570
rect 8740 173270 8800 173570
rect 9100 173270 9160 173570
rect 9460 173270 9520 173570
rect 9820 173270 9880 173570
rect 10180 173270 10240 173570
rect 10540 173270 10600 173570
rect 10900 173270 10960 173570
rect 11260 173270 11320 173570
rect 11620 173270 11680 173570
rect 11980 173270 12000 173570
rect 8000 173210 12000 173270
rect 8000 172910 8080 173210
rect 8380 172910 8440 173210
rect 8740 172910 8800 173210
rect 9100 172910 9160 173210
rect 9460 172910 9520 173210
rect 9820 172910 9880 173210
rect 10180 172910 10240 173210
rect 10540 172910 10600 173210
rect 10900 172910 10960 173210
rect 11260 172910 11320 173210
rect 11620 172910 11680 173210
rect 11980 172910 12000 173210
rect 8000 172000 12000 172910
rect 109388 16020 112268 423040
rect 109388 15580 110600 16020
rect 111040 15580 112268 16020
rect 109388 15520 112268 15580
rect 109388 15080 110600 15520
rect 111040 15080 112268 15520
rect 109388 15020 112268 15080
rect 109388 14580 110600 15020
rect 111040 14580 112268 15020
rect 109388 14520 112268 14580
rect 109388 14080 110600 14520
rect 111040 14080 112268 14520
rect 109388 14020 112268 14080
rect 109388 13580 110600 14020
rect 111040 13580 112268 14020
rect 109388 13520 112268 13580
rect 109388 13080 110600 13520
rect 111040 13080 112268 13520
rect 109388 13020 112268 13080
rect 109388 12580 110600 13020
rect 111040 12580 112268 13020
rect 109388 12520 112268 12580
rect 109388 12080 110600 12520
rect 111040 12080 112268 12520
rect 109388 12000 112268 12080
rect 113706 16020 116408 423882
rect 113706 15580 114810 16020
rect 115250 15580 116408 16020
rect 113706 15520 116408 15580
rect 113706 15080 114810 15520
rect 115250 15080 116408 15520
rect 113706 15020 116408 15080
rect 113706 14580 114810 15020
rect 115250 14580 116408 15020
rect 113706 14520 116408 14580
rect 113706 14080 114810 14520
rect 115250 14080 116408 14520
rect 113706 14020 116408 14080
rect 113706 13580 114810 14020
rect 115250 13580 116408 14020
rect 113706 13520 116408 13580
rect 113706 13080 114810 13520
rect 115250 13080 116408 13520
rect 113706 13020 116408 13080
rect 113706 12580 114810 13020
rect 115250 12580 116408 13020
rect 113706 12520 116408 12580
rect 113706 12080 114810 12520
rect 115250 12080 116408 12520
rect 113706 12000 116408 12080
rect 118266 16020 120678 420078
rect 118266 15580 119240 16020
rect 119680 15580 120678 16020
rect 118266 15520 120678 15580
rect 118266 15080 119240 15520
rect 119680 15080 120678 15520
rect 118266 15020 120678 15080
rect 118266 14580 119240 15020
rect 119680 14580 120678 15020
rect 118266 14520 120678 14580
rect 118266 14080 119240 14520
rect 119680 14080 120678 14520
rect 118266 14020 120678 14080
rect 118266 13580 119240 14020
rect 119680 13580 120678 14020
rect 118266 13520 120678 13580
rect 118266 13080 119240 13520
rect 119680 13080 120678 13520
rect 118266 13020 120678 13080
rect 118266 12580 119240 13020
rect 119680 12580 120678 13020
rect 118266 12520 120678 12580
rect 118266 12080 119240 12520
rect 119680 12080 120678 12520
rect 118266 12000 120678 12080
rect 122404 16020 125264 417212
rect 122404 15580 123600 16020
rect 124040 15580 125264 16020
rect 122404 15520 125264 15580
rect 122404 15080 123600 15520
rect 124040 15080 125264 15520
rect 122404 15020 125264 15080
rect 122404 14580 123600 15020
rect 124040 14580 125264 15020
rect 122404 14520 125264 14580
rect 122404 14080 123600 14520
rect 124040 14080 125264 14520
rect 122404 14020 125264 14080
rect 122404 13580 123600 14020
rect 124040 13580 125264 14020
rect 122404 13520 125264 13580
rect 122404 13080 123600 13520
rect 124040 13080 125264 13520
rect 122404 13020 125264 13080
rect 122404 12580 123600 13020
rect 124040 12580 125264 13020
rect 122404 12520 125264 12580
rect 122404 12080 123600 12520
rect 124040 12080 125264 12520
rect 122404 12000 125264 12080
rect 126932 16020 129668 413392
rect 131176 35150 134144 409064
rect 131176 34550 131200 35150
rect 131800 34550 131960 35150
rect 132560 34550 132740 35150
rect 133340 34550 133500 35150
rect 134100 34550 134144 35150
rect 131176 34450 134144 34550
rect 126932 15580 128080 16020
rect 128520 15580 129668 16020
rect 126932 15520 129668 15580
rect 126932 15080 128080 15520
rect 128520 15080 129668 15520
rect 126932 15020 129668 15080
rect 126932 14580 128080 15020
rect 128520 14580 129668 15020
rect 126932 14520 129668 14580
rect 126932 14080 128080 14520
rect 128520 14080 129668 14520
rect 126932 14020 129668 14080
rect 126932 13580 128080 14020
rect 128520 13580 129668 14020
rect 126932 13520 129668 13580
rect 126932 13080 128080 13520
rect 128520 13080 129668 13520
rect 126932 13020 129668 13080
rect 126932 12580 128080 13020
rect 128520 12580 129668 13020
rect 126932 12520 129668 12580
rect 126932 12080 128080 12520
rect 128520 12080 129668 12520
rect 126932 12000 129668 12080
rect 135890 14646 138534 406444
rect 156892 371880 159750 384150
rect 156892 371580 156900 371880
rect 157200 371580 157260 371880
rect 157560 371580 157620 371880
rect 157920 371580 157980 371880
rect 158280 371580 158340 371880
rect 158640 371580 158700 371880
rect 159000 371580 159060 371880
rect 159360 371580 159420 371880
rect 159720 371580 159750 371880
rect 156892 371520 159750 371580
rect 156892 371220 156900 371520
rect 157200 371220 157260 371520
rect 157560 371220 157620 371520
rect 157920 371220 157980 371520
rect 158280 371220 158340 371520
rect 158640 371220 158700 371520
rect 159000 371220 159060 371520
rect 159360 371220 159420 371520
rect 159720 371220 159750 371520
rect 156892 371160 159750 371220
rect 156892 370860 156900 371160
rect 157200 370860 157260 371160
rect 157560 370860 157620 371160
rect 157920 370860 157980 371160
rect 158280 370860 158340 371160
rect 158640 370860 158700 371160
rect 159000 370860 159060 371160
rect 159360 370860 159420 371160
rect 159720 370860 159750 371160
rect 156892 370800 159750 370860
rect 156892 370500 156900 370800
rect 157200 370500 157260 370800
rect 157560 370500 157620 370800
rect 157920 370500 157980 370800
rect 158280 370500 158340 370800
rect 158640 370500 158700 370800
rect 159000 370500 159060 370800
rect 159360 370500 159420 370800
rect 159720 370500 159750 370800
rect 156892 370440 159750 370500
rect 156892 370140 156900 370440
rect 157200 370140 157260 370440
rect 157560 370140 157620 370440
rect 157920 370140 157980 370440
rect 158280 370140 158340 370440
rect 158640 370140 158700 370440
rect 159000 370140 159060 370440
rect 159360 370140 159420 370440
rect 159720 370140 159750 370440
rect 156892 370080 159750 370140
rect 156892 369780 156900 370080
rect 157200 369780 157260 370080
rect 157560 369780 157620 370080
rect 157920 369780 157980 370080
rect 158280 369780 158340 370080
rect 158640 369780 158700 370080
rect 159000 369780 159060 370080
rect 159360 369780 159420 370080
rect 159720 369780 159750 370080
rect 156892 369760 159750 369780
rect 232714 366414 235572 384411
rect 232714 366114 232722 366414
rect 233022 366114 233082 366414
rect 233382 366114 233442 366414
rect 233742 366114 233802 366414
rect 234102 366114 234162 366414
rect 234462 366114 234522 366414
rect 234822 366114 234882 366414
rect 235182 366114 235242 366414
rect 235542 366114 235572 366414
rect 232714 366054 235572 366114
rect 232714 365754 232722 366054
rect 233022 365754 233082 366054
rect 233382 365754 233442 366054
rect 233742 365754 233802 366054
rect 234102 365754 234162 366054
rect 234462 365754 234522 366054
rect 234822 365754 234882 366054
rect 235182 365754 235242 366054
rect 235542 365754 235572 366054
rect 232714 365694 235572 365754
rect 232714 365394 232722 365694
rect 233022 365394 233082 365694
rect 233382 365394 233442 365694
rect 233742 365394 233802 365694
rect 234102 365394 234162 365694
rect 234462 365394 234522 365694
rect 234822 365394 234882 365694
rect 235182 365394 235242 365694
rect 235542 365394 235572 365694
rect 232714 365334 235572 365394
rect 232714 365034 232722 365334
rect 233022 365034 233082 365334
rect 233382 365034 233442 365334
rect 233742 365034 233802 365334
rect 234102 365034 234162 365334
rect 234462 365034 234522 365334
rect 234822 365034 234882 365334
rect 235182 365034 235242 365334
rect 235542 365034 235572 365334
rect 232714 364974 235572 365034
rect 232714 364674 232722 364974
rect 233022 364674 233082 364974
rect 233382 364674 233442 364974
rect 233742 364674 233802 364974
rect 234102 364674 234162 364974
rect 234462 364674 234522 364974
rect 234822 364674 234882 364974
rect 235182 364674 235242 364974
rect 235542 364674 235572 364974
rect 232714 364614 235572 364674
rect 232714 364314 232722 364614
rect 233022 364314 233082 364614
rect 233382 364314 233442 364614
rect 233742 364314 233802 364614
rect 234102 364314 234162 364614
rect 234462 364314 234522 364614
rect 234822 364314 234882 364614
rect 235182 364314 235242 364614
rect 235542 364314 235572 364614
rect 232714 364280 235572 364314
rect 310508 360188 313366 388534
rect 310508 359888 310516 360188
rect 310816 359888 310876 360188
rect 311176 359888 311236 360188
rect 311536 359888 311596 360188
rect 311896 359888 311956 360188
rect 312256 359888 312316 360188
rect 312616 359888 312676 360188
rect 312976 359888 313036 360188
rect 313336 359888 313366 360188
rect 310508 359828 313366 359888
rect 310508 359528 310516 359828
rect 310816 359528 310876 359828
rect 311176 359528 311236 359828
rect 311536 359528 311596 359828
rect 311896 359528 311956 359828
rect 312256 359528 312316 359828
rect 312616 359528 312676 359828
rect 312976 359528 313036 359828
rect 313336 359528 313366 359828
rect 310508 359468 313366 359528
rect 310508 359168 310516 359468
rect 310816 359168 310876 359468
rect 311176 359168 311236 359468
rect 311536 359168 311596 359468
rect 311896 359168 311956 359468
rect 312256 359168 312316 359468
rect 312616 359168 312676 359468
rect 312976 359168 313036 359468
rect 313336 359168 313366 359468
rect 310508 359108 313366 359168
rect 310508 358808 310516 359108
rect 310816 358808 310876 359108
rect 311176 358808 311236 359108
rect 311536 358808 311596 359108
rect 311896 358808 311956 359108
rect 312256 358808 312316 359108
rect 312616 358808 312676 359108
rect 312976 358808 313036 359108
rect 313336 358808 313366 359108
rect 310508 358748 313366 358808
rect 310508 358448 310516 358748
rect 310816 358448 310876 358748
rect 311176 358448 311236 358748
rect 311536 358448 311596 358748
rect 311896 358448 311956 358748
rect 312256 358448 312316 358748
rect 312616 358448 312676 358748
rect 312976 358448 313036 358748
rect 313336 358448 313366 358748
rect 310508 358388 313366 358448
rect 310508 358088 310516 358388
rect 310816 358088 310876 358388
rect 311176 358088 311236 358388
rect 311536 358088 311596 358388
rect 311896 358088 311956 358388
rect 312256 358088 312316 358388
rect 312616 358088 312676 358388
rect 312976 358088 313036 358388
rect 313336 358088 313366 358388
rect 310508 358020 313366 358088
rect 135890 14520 145038 14646
rect 135890 14080 144562 14520
rect 145002 14080 145038 14520
rect 135890 14020 145038 14080
rect 135890 13580 144562 14020
rect 145002 13580 145038 14020
rect 135890 13520 145038 13580
rect 135890 13080 144562 13520
rect 145002 13080 145038 13520
rect 135890 13020 145038 13080
rect 135890 12580 144562 13020
rect 145002 12580 145038 13020
rect 135890 12520 145038 12580
rect 135890 12080 144562 12520
rect 145002 12080 145038 12520
rect 135890 12002 145038 12080
rect 144522 12000 145012 12002
<< via4 >>
rect 16200 582600 23800 582800
rect 16200 575400 16400 582600
rect 16400 575400 23600 582600
rect 23600 575400 23800 582600
rect 16200 575200 23800 575400
rect 16200 558200 23800 565800
rect 109480 424640 109780 424940
rect 109880 424640 110180 424940
rect 110280 424640 110580 424940
rect 110680 424640 110980 424940
rect 111080 424640 111380 424940
rect 111480 424640 111780 424940
rect 111880 424640 112180 424940
rect 109480 424240 109780 424540
rect 109880 424240 110180 424540
rect 110280 424240 110580 424540
rect 110680 424240 110980 424540
rect 111080 424240 111380 424540
rect 111480 424240 111780 424540
rect 111880 424240 112180 424540
rect 109480 423840 109780 424140
rect 109880 423840 110180 424140
rect 110280 423840 110580 424140
rect 110680 423840 110980 424140
rect 111080 423840 111380 424140
rect 111480 423840 111780 424140
rect 111880 423840 112180 424140
rect 109480 423440 109780 423740
rect 109880 423440 110180 423740
rect 110280 423440 110580 423740
rect 110680 423440 110980 423740
rect 111080 423440 111380 423740
rect 111480 423440 111780 423740
rect 111880 423440 112180 423740
rect 109480 423040 109780 423340
rect 109880 423040 110180 423340
rect 110280 423040 110580 423340
rect 110680 423040 110980 423340
rect 111080 423040 111380 423340
rect 111480 423040 111780 423340
rect 111880 423040 112180 423340
rect 31028 400264 31628 400274
rect 31028 399704 31048 400264
rect 31048 399704 31608 400264
rect 31608 399704 31628 400264
rect 31028 399674 31628 399704
rect 31728 400264 32328 400274
rect 31728 399704 31748 400264
rect 31748 399704 32308 400264
rect 32308 399704 32328 400264
rect 31728 399674 32328 399704
rect 32428 400264 33028 400274
rect 32428 399704 32448 400264
rect 32448 399704 33008 400264
rect 33008 399704 33028 400264
rect 32428 399674 33028 399704
rect 33128 400264 33728 400274
rect 33128 399704 33148 400264
rect 33148 399704 33708 400264
rect 33708 399704 33728 400264
rect 33128 399674 33728 399704
rect 31028 399564 31628 399574
rect 31028 399004 31048 399564
rect 31048 399004 31608 399564
rect 31608 399004 31628 399564
rect 31028 398974 31628 399004
rect 31728 399564 32328 399574
rect 31728 399004 31748 399564
rect 31748 399004 32308 399564
rect 32308 399004 32328 399564
rect 31728 398974 32328 399004
rect 32428 399564 33028 399574
rect 32428 399004 32448 399564
rect 32448 399004 33008 399564
rect 33008 399004 33028 399564
rect 32428 398974 33028 399004
rect 33128 399564 33728 399574
rect 33128 399004 33148 399564
rect 33148 399004 33708 399564
rect 33708 399004 33728 399564
rect 33128 398974 33728 399004
rect 31028 398864 31628 398874
rect 31028 398304 31048 398864
rect 31048 398304 31608 398864
rect 31608 398304 31628 398864
rect 31028 398274 31628 398304
rect 31728 398864 32328 398874
rect 31728 398304 31748 398864
rect 31748 398304 32308 398864
rect 32308 398304 32328 398864
rect 31728 398274 32328 398304
rect 32428 398864 33028 398874
rect 32428 398304 32448 398864
rect 32448 398304 33008 398864
rect 33008 398304 33028 398864
rect 32428 398274 33028 398304
rect 33128 398864 33728 398874
rect 33128 398304 33148 398864
rect 33148 398304 33708 398864
rect 33708 398304 33728 398864
rect 33128 398274 33728 398304
rect 31000 396778 31600 396788
rect 31000 396218 31020 396778
rect 31020 396218 31580 396778
rect 31580 396218 31600 396778
rect 31000 396188 31600 396218
rect 31700 396778 32300 396788
rect 31700 396218 31720 396778
rect 31720 396218 32280 396778
rect 32280 396218 32300 396778
rect 31700 396188 32300 396218
rect 32400 396778 33000 396788
rect 32400 396218 32420 396778
rect 32420 396218 32980 396778
rect 32980 396218 33000 396778
rect 32400 396188 33000 396218
rect 33100 396778 33700 396788
rect 33100 396218 33120 396778
rect 33120 396218 33680 396778
rect 33680 396218 33700 396778
rect 33100 396188 33700 396218
rect 31000 396078 31600 396088
rect 31000 395518 31020 396078
rect 31020 395518 31580 396078
rect 31580 395518 31600 396078
rect 31000 395488 31600 395518
rect 31700 396078 32300 396088
rect 31700 395518 31720 396078
rect 31720 395518 32280 396078
rect 32280 395518 32300 396078
rect 31700 395488 32300 395518
rect 32400 396078 33000 396088
rect 32400 395518 32420 396078
rect 32420 395518 32980 396078
rect 32980 395518 33000 396078
rect 32400 395488 33000 395518
rect 33100 396078 33700 396088
rect 33100 395518 33120 396078
rect 33120 395518 33680 396078
rect 33680 395518 33700 396078
rect 33100 395488 33700 395518
rect 31000 395378 31600 395388
rect 31000 394818 31020 395378
rect 31020 394818 31580 395378
rect 31580 394818 31600 395378
rect 31000 394788 31600 394818
rect 31700 395378 32300 395388
rect 31700 394818 31720 395378
rect 31720 394818 32280 395378
rect 32280 394818 32300 395378
rect 31700 394788 32300 394818
rect 32400 395378 33000 395388
rect 32400 394818 32420 395378
rect 32420 394818 32980 395378
rect 32980 394818 33000 395378
rect 32400 394788 33000 394818
rect 33100 395378 33700 395388
rect 33100 394818 33120 395378
rect 33120 394818 33680 395378
rect 33680 394818 33700 395378
rect 33100 394788 33700 394818
rect 31068 393138 31668 393148
rect 31068 392578 31088 393138
rect 31088 392578 31648 393138
rect 31648 392578 31668 393138
rect 31068 392548 31668 392578
rect 31768 393138 32368 393148
rect 31768 392578 31788 393138
rect 31788 392578 32348 393138
rect 32348 392578 32368 393138
rect 31768 392548 32368 392578
rect 32468 393138 33068 393148
rect 32468 392578 32488 393138
rect 32488 392578 33048 393138
rect 33048 392578 33068 393138
rect 32468 392548 33068 392578
rect 33168 393138 33768 393148
rect 33168 392578 33188 393138
rect 33188 392578 33748 393138
rect 33748 392578 33768 393138
rect 33168 392548 33768 392578
rect 31068 392438 31668 392448
rect 31068 391878 31088 392438
rect 31088 391878 31648 392438
rect 31648 391878 31668 392438
rect 31068 391848 31668 391878
rect 31768 392438 32368 392448
rect 31768 391878 31788 392438
rect 31788 391878 32348 392438
rect 32348 391878 32368 392438
rect 31768 391848 32368 391878
rect 32468 392438 33068 392448
rect 32468 391878 32488 392438
rect 32488 391878 33048 392438
rect 33048 391878 33068 392438
rect 32468 391848 33068 391878
rect 33168 392438 33768 392448
rect 33168 391878 33188 392438
rect 33188 391878 33748 392438
rect 33748 391878 33768 392438
rect 33168 391848 33768 391878
rect 31068 391738 31668 391748
rect 31068 391178 31088 391738
rect 31088 391178 31648 391738
rect 31648 391178 31668 391738
rect 31068 391148 31668 391178
rect 31768 391738 32368 391748
rect 31768 391178 31788 391738
rect 31788 391178 32348 391738
rect 32348 391178 32368 391738
rect 31768 391148 32368 391178
rect 32468 391738 33068 391748
rect 32468 391178 32488 391738
rect 32488 391178 33048 391738
rect 33048 391178 33068 391738
rect 32468 391148 33068 391178
rect 33168 391738 33768 391748
rect 33168 391178 33188 391738
rect 33188 391178 33748 391738
rect 33748 391178 33768 391738
rect 33168 391148 33768 391178
rect 31068 389034 31668 389044
rect 31068 388474 31088 389034
rect 31088 388474 31648 389034
rect 31648 388474 31668 389034
rect 31068 388444 31668 388474
rect 31768 389034 32368 389044
rect 31768 388474 31788 389034
rect 31788 388474 32348 389034
rect 32348 388474 32368 389034
rect 31768 388444 32368 388474
rect 32468 389034 33068 389044
rect 32468 388474 32488 389034
rect 32488 388474 33048 389034
rect 33048 388474 33068 389034
rect 32468 388444 33068 388474
rect 33168 389034 33768 389044
rect 33168 388474 33188 389034
rect 33188 388474 33748 389034
rect 33748 388474 33768 389034
rect 33168 388444 33768 388474
rect 31068 388334 31668 388344
rect 31068 387774 31088 388334
rect 31088 387774 31648 388334
rect 31648 387774 31668 388334
rect 31068 387744 31668 387774
rect 31768 388334 32368 388344
rect 31768 387774 31788 388334
rect 31788 387774 32348 388334
rect 32348 387774 32368 388334
rect 31768 387744 32368 387774
rect 32468 388334 33068 388344
rect 32468 387774 32488 388334
rect 32488 387774 33048 388334
rect 33048 387774 33068 388334
rect 32468 387744 33068 387774
rect 33168 388334 33768 388344
rect 33168 387774 33188 388334
rect 33188 387774 33748 388334
rect 33748 387774 33768 388334
rect 33168 387744 33768 387774
rect 31068 387634 31668 387644
rect 31068 387074 31088 387634
rect 31088 387074 31648 387634
rect 31648 387074 31668 387634
rect 31068 387044 31668 387074
rect 31768 387634 32368 387644
rect 31768 387074 31788 387634
rect 31788 387074 32348 387634
rect 32348 387074 32368 387634
rect 31768 387044 32368 387074
rect 32468 387634 33068 387644
rect 32468 387074 32488 387634
rect 32488 387074 33048 387634
rect 33048 387074 33068 387634
rect 32468 387044 33068 387074
rect 33168 387634 33768 387644
rect 33168 387074 33188 387634
rect 33188 387074 33748 387634
rect 33748 387074 33768 387634
rect 33168 387044 33768 387074
rect 31200 385590 31800 385600
rect 31200 385030 31220 385590
rect 31220 385030 31780 385590
rect 31780 385030 31800 385590
rect 31200 385000 31800 385030
rect 31900 385590 32500 385600
rect 31900 385030 31920 385590
rect 31920 385030 32480 385590
rect 32480 385030 32500 385590
rect 31900 385000 32500 385030
rect 32600 385590 33200 385600
rect 32600 385030 32620 385590
rect 32620 385030 33180 385590
rect 33180 385030 33200 385590
rect 32600 385000 33200 385030
rect 33300 385590 33900 385600
rect 33300 385030 33320 385590
rect 33320 385030 33880 385590
rect 33880 385030 33900 385590
rect 33300 385000 33900 385030
rect 31200 384890 31800 384900
rect 31200 384330 31220 384890
rect 31220 384330 31780 384890
rect 31780 384330 31800 384890
rect 31200 384300 31800 384330
rect 31900 384890 32500 384900
rect 31900 384330 31920 384890
rect 31920 384330 32480 384890
rect 32480 384330 32500 384890
rect 31900 384300 32500 384330
rect 32600 384890 33200 384900
rect 32600 384330 32620 384890
rect 32620 384330 33180 384890
rect 33180 384330 33200 384890
rect 32600 384300 33200 384330
rect 33300 384890 33900 384900
rect 33300 384330 33320 384890
rect 33320 384330 33880 384890
rect 33880 384330 33900 384890
rect 33300 384300 33900 384330
rect 31200 384190 31800 384200
rect 31200 383630 31220 384190
rect 31220 383630 31780 384190
rect 31780 383630 31800 384190
rect 31200 383600 31800 383630
rect 31900 384190 32500 384200
rect 31900 383630 31920 384190
rect 31920 383630 32480 384190
rect 32480 383630 32500 384190
rect 31900 383600 32500 383630
rect 32600 384190 33200 384200
rect 32600 383630 32620 384190
rect 32620 383630 33180 384190
rect 33180 383630 33200 384190
rect 32600 383600 33200 383630
rect 33300 384190 33900 384200
rect 33300 383630 33320 384190
rect 33320 383630 33880 384190
rect 33880 383630 33900 384190
rect 33300 383600 33900 383630
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 16000 582800 24000 583000
rect 16000 575200 16200 582800
rect 23800 575200 24000 582800
rect 16000 575000 24000 575200
rect 16000 565800 24000 566000
rect 16000 558200 16200 565800
rect 23800 558200 24000 565800
rect 16000 558000 24000 558200
rect 109388 424940 112268 425000
rect 109388 424640 109480 424940
rect 109780 424640 109880 424940
rect 110180 424640 110280 424940
rect 110580 424640 110680 424940
rect 110980 424640 111080 424940
rect 111380 424640 111480 424940
rect 111780 424640 111880 424940
rect 112180 424640 112268 424940
rect 109388 424540 112268 424640
rect 109388 424240 109480 424540
rect 109780 424240 109880 424540
rect 110180 424240 110280 424540
rect 110580 424240 110680 424540
rect 110980 424240 111080 424540
rect 111380 424240 111480 424540
rect 111780 424240 111880 424540
rect 112180 424240 112268 424540
rect 109388 424140 112268 424240
rect 109388 423840 109480 424140
rect 109780 423840 109880 424140
rect 110180 423840 110280 424140
rect 110580 423840 110680 424140
rect 110980 423840 111080 424140
rect 111380 423840 111480 424140
rect 111780 423840 111880 424140
rect 112180 423840 112268 424140
rect 109388 423740 112268 423840
rect 109388 423440 109480 423740
rect 109780 423440 109880 423740
rect 110180 423440 110280 423740
rect 110580 423440 110680 423740
rect 110980 423440 111080 423740
rect 111380 423440 111480 423740
rect 111780 423440 111880 423740
rect 112180 423440 112268 423740
rect 109388 423340 112268 423440
rect 109388 423040 109480 423340
rect 109780 423040 109880 423340
rect 110180 423040 110280 423340
rect 110580 423040 110680 423340
rect 110980 423040 111080 423340
rect 111380 423040 111480 423340
rect 111780 423040 111880 423340
rect 112180 423040 112268 423340
rect 109388 422980 112268 423040
rect 30988 400274 33768 400314
rect 30988 399674 31028 400274
rect 31628 399674 31728 400274
rect 32328 399674 32428 400274
rect 33028 399674 33128 400274
rect 33728 399674 33768 400274
rect 30988 399574 33768 399674
rect 30988 398974 31028 399574
rect 31628 398974 31728 399574
rect 32328 398974 32428 399574
rect 33028 398974 33128 399574
rect 33728 398974 33768 399574
rect 30988 398874 33768 398974
rect 30988 398274 31028 398874
rect 31628 398274 31728 398874
rect 32328 398274 32428 398874
rect 33028 398274 33128 398874
rect 33728 398274 33768 398874
rect 30988 398244 33768 398274
rect 30960 396788 33740 396828
rect 30960 396188 31000 396788
rect 31600 396188 31700 396788
rect 32300 396188 32400 396788
rect 33000 396188 33100 396788
rect 33700 396188 33740 396788
rect 30960 396088 33740 396188
rect 30960 395488 31000 396088
rect 31600 395488 31700 396088
rect 32300 395488 32400 396088
rect 33000 395488 33100 396088
rect 33700 395488 33740 396088
rect 30960 395388 33740 395488
rect 30960 394788 31000 395388
rect 31600 394788 31700 395388
rect 32300 394788 32400 395388
rect 33000 394788 33100 395388
rect 33700 394788 33740 395388
rect 30960 394758 33740 394788
rect 31028 393148 33808 393188
rect 31028 392548 31068 393148
rect 31668 392548 31768 393148
rect 32368 392548 32468 393148
rect 33068 392548 33168 393148
rect 33768 392548 33808 393148
rect 31028 392448 33808 392548
rect 31028 391848 31068 392448
rect 31668 391848 31768 392448
rect 32368 391848 32468 392448
rect 33068 391848 33168 392448
rect 33768 391848 33808 392448
rect 31028 391748 33808 391848
rect 31028 391148 31068 391748
rect 31668 391148 31768 391748
rect 32368 391148 32468 391748
rect 33068 391148 33168 391748
rect 33768 391148 33808 391748
rect 31028 391118 33808 391148
rect 31028 389044 33808 389084
rect 31028 388444 31068 389044
rect 31668 388444 31768 389044
rect 32368 388444 32468 389044
rect 33068 388444 33168 389044
rect 33768 388444 33808 389044
rect 31028 388344 33808 388444
rect 31028 387744 31068 388344
rect 31668 387744 31768 388344
rect 32368 387744 32468 388344
rect 33068 387744 33168 388344
rect 33768 387744 33808 388344
rect 31028 387644 33808 387744
rect 31028 387044 31068 387644
rect 31668 387044 31768 387644
rect 32368 387044 32468 387644
rect 33068 387044 33168 387644
rect 33768 387044 33808 387644
rect 31028 387014 33808 387044
rect 31160 385600 33940 385640
rect 31160 385000 31200 385600
rect 31800 385000 31900 385600
rect 32500 385000 32600 385600
rect 33200 385000 33300 385600
rect 33900 385000 33940 385600
rect 31160 384900 33940 385000
rect 31160 384300 31200 384900
rect 31800 384300 31900 384900
rect 32500 384300 32600 384900
rect 33200 384300 33300 384900
rect 33900 384300 33940 384900
rect 31160 384200 33940 384300
rect 31160 383600 31200 384200
rect 31800 383600 31900 384200
rect 32500 383600 32600 384200
rect 33200 383600 33300 384200
rect 33900 383600 33940 384200
rect 31160 383570 33940 383600
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect 586000 586000 588000 588000
rect 586000 496000 588000 498000
rect 586000 452000 588000 454000
rect 586000 406000 588000 408000
rect -100 -100 584100 0
use MulColROs  MulColROs_0 ../user_prj/MulColRO/mag
timestamp 1698914393
transform 1 0 -40398 0 1 -219150
box 62168 599934 367990 811050
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
