magic
tech sky130A
magscale 1 2
timestamp 1699164000
<< metal4 >>
rect -3000 8000 3000 8057
rect -3000 -8057 3000 -8000
<< rmetal4 >>
rect -3000 -8000 3000 8000
<< properties >>
string gencell sky130_fd_pr__res_generic_m4
string library sky130
string parameters w 30.0 l 80.0 m 1 nx 1 wmin 0.30 lmin 0.30 rho 0.047 val 125.333m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
