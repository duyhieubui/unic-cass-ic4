magic
tech sky130A
magscale 1 2
timestamp 1699297357
<< isosubstrate >>
rect 385684 591732 438400 634000
rect 463604 542910 544568 544424
rect 50782 326818 356604 537934
rect 463604 506200 547380 542910
rect 463604 500600 529000 506200
rect 540800 500600 547380 506200
rect 463604 495830 547380 500600
rect 469516 492874 547380 495830
<< metal2 >>
rect 381271 616766 387143 618225
rect 381271 571010 382730 616766
rect 384041 614573 386359 614891
rect 384041 573410 384359 614573
rect 385641 612519 386359 612837
rect 385642 575410 385958 612519
rect 385600 575400 386000 575410
rect 385600 574990 386000 575000
rect 384000 573400 384400 573410
rect 384000 572990 384400 573000
rect 381000 571000 383000 571010
rect 381000 568990 383000 569000
rect 570300 319900 570900 319910
rect 118620 16000 119020 16010
rect 122830 16000 123230 16010
rect 127260 16000 127660 16010
rect 131620 16000 132020 16010
rect 136100 16000 136500 16010
rect 119020 15600 119030 16000
rect 118620 15500 119030 15600
rect 119020 15100 119030 15500
rect 118620 15000 119030 15100
rect 119020 14600 119030 15000
rect 118620 14500 119030 14600
rect 119020 14100 119030 14500
rect 118620 14000 119030 14100
rect 119020 13600 119030 14000
rect 118620 13500 119030 13600
rect 119020 13100 119030 13500
rect 118620 13000 119030 13100
rect 119020 12600 119030 13000
rect 118620 12500 119030 12600
rect 119020 12100 119030 12500
rect 118620 2401 119030 12100
rect 123230 15600 123250 16000
rect 122830 15500 123250 15600
rect 123230 15100 123250 15500
rect 122830 15000 123250 15100
rect 123230 14600 123250 15000
rect 122830 14500 123250 14600
rect 123230 14100 123250 14500
rect 122830 14000 123250 14100
rect 123230 13600 123250 14000
rect 122830 13500 123250 13600
rect 123230 13100 123250 13500
rect 122830 13000 123250 13100
rect 123230 12600 123250 13000
rect 122830 12500 123250 12600
rect 123230 12100 123250 12500
rect 122830 4409 123250 12100
rect 127660 15600 127670 16000
rect 127260 15500 127670 15600
rect 127660 15100 127670 15500
rect 127260 15000 127670 15100
rect 127660 14600 127670 15000
rect 127260 14500 127670 14600
rect 127660 14100 127670 14500
rect 127260 14000 127670 14100
rect 127660 13600 127670 14000
rect 127260 13500 127670 13600
rect 127660 13100 127670 13500
rect 127260 13000 127670 13100
rect 127660 12600 127670 13000
rect 127260 12500 127670 12600
rect 127660 12100 127670 12500
rect 127260 6399 127670 12100
rect 132020 15600 132030 16000
rect 131620 15500 132030 15600
rect 132020 15100 132030 15500
rect 131620 15000 132030 15100
rect 132020 14600 132030 15000
rect 131620 14500 132030 14600
rect 132020 14100 132030 14500
rect 131620 14000 132030 14100
rect 132020 13600 132030 14000
rect 131620 13500 132030 13600
rect 132020 13100 132030 13500
rect 131620 13000 132030 13100
rect 132020 12600 132030 13000
rect 131620 12500 132030 12600
rect 132020 12100 132030 12500
rect 131620 8400 132030 12100
rect 136500 15600 136510 16000
rect 136100 15500 136510 15600
rect 136500 15100 136510 15500
rect 136100 15000 136510 15100
rect 136500 14600 136510 15000
rect 136100 14500 136510 14600
rect 136500 14100 136510 14500
rect 136100 14000 136510 14100
rect 136500 13600 136510 14000
rect 136100 13500 136510 13600
rect 136500 13100 136510 13500
rect 136100 13000 136510 13100
rect 136500 12600 136510 13000
rect 136100 12500 136510 12600
rect 136500 12100 136510 12500
rect 136100 10400 136510 12100
rect 144582 14500 144982 14536
rect 144582 14000 144982 14100
rect 144582 13500 144982 13600
rect 144582 13000 144982 13100
rect 144582 12500 144982 12600
rect 136100 10000 141432 10400
rect 131620 8000 137882 8400
rect 127260 6000 134340 6399
rect 122830 4009 130800 4409
rect 122830 4000 127252 4009
rect 128000 4000 130800 4009
rect 118620 2000 127250 2401
rect 126850 790 127250 2000
rect 126860 780 127250 790
rect 126870 770 127240 780
rect 126880 760 127230 770
rect 126890 750 127220 760
rect 126900 740 127210 750
rect 130390 740 130800 4000
rect 133940 740 134340 6000
rect 137482 740 137882 8000
rect 141032 780 141432 10000
rect 144582 810 144982 12100
rect 570300 7400 570900 319300
rect 570300 5400 570900 6400
rect 144592 800 144982 810
rect 566500 4800 570900 5400
rect 571900 275500 572500 275510
rect 571900 7400 572500 274900
rect 566500 800 567100 4800
rect 571900 3800 572500 6400
rect 570000 3200 572500 3800
rect 573500 95400 574100 95410
rect 573500 7400 574100 94800
rect 570000 800 570600 3200
rect 573500 800 574100 6400
rect 575100 50800 575700 50810
rect 575100 7400 575700 50200
rect 575100 3800 575700 6400
rect 575100 3200 577700 3800
rect 577100 800 577700 3200
rect 144602 790 144972 800
rect 144612 780 144962 790
rect 141042 770 141432 780
rect 144622 770 144952 780
rect 141052 760 141422 770
rect 144632 760 144942 770
rect 141062 750 141412 760
rect 144642 750 144932 760
rect 141072 740 141402 750
rect 144652 740 144922 750
rect 126910 730 127200 740
rect 130400 730 130800 740
rect 133950 730 134340 740
rect 137492 730 137882 740
rect 141082 730 141392 740
rect 144662 730 144912 740
rect 126920 720 127190 730
rect 130410 720 130790 730
rect 133960 720 134330 730
rect 137502 720 137872 730
rect 141092 720 141382 730
rect 144672 720 144902 730
rect 126930 710 127180 720
rect 130420 710 130780 720
rect 133970 710 134320 720
rect 137512 710 137862 720
rect 141102 710 141372 720
rect 144682 710 144892 720
rect 126940 700 127170 710
rect 130430 700 130770 710
rect 133980 700 134310 710
rect 137522 700 137852 710
rect 141112 700 141362 710
rect 144692 700 144882 710
rect 126950 690 127160 700
rect 130440 690 130760 700
rect 133990 690 134300 700
rect 137532 690 137842 700
rect 141122 690 141352 700
rect 144702 690 144872 700
rect 126960 680 127150 690
rect 130450 680 130750 690
rect 134000 680 134290 690
rect 137542 680 137832 690
rect 141132 680 141342 690
rect 144712 680 144862 690
rect 126970 670 127140 680
rect 130460 670 130740 680
rect 134010 670 134280 680
rect 137552 670 137822 680
rect 141142 670 141332 680
rect 144722 670 144852 680
rect 126980 660 127130 670
rect 130470 660 130730 670
rect 134020 660 134270 670
rect 137562 660 137812 670
rect 141152 660 141322 670
rect 126990 650 127120 660
rect 130480 650 130720 660
rect 134030 650 134260 660
rect 137572 650 137802 660
rect 141162 650 141312 660
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 650
rect 130490 640 130710 650
rect 134040 640 134250 650
rect 137582 640 137792 650
rect 141172 640 141302 650
rect 130500 630 130700 640
rect 134050 630 134240 640
rect 137592 630 137782 640
rect 130510 620 130690 630
rect 134060 620 134230 630
rect 137602 620 137772 630
rect 130520 610 130680 620
rect 134070 610 134220 620
rect 137612 610 137762 620
rect 130530 600 130670 610
rect 134080 600 134210 610
rect 137622 600 137752 610
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 600
rect 131726 -800 131838 480
rect 132908 -800 133020 600
rect 134090 -800 134202 600
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 600
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 640
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 670
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 800
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 800
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 800
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 800
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< rmetal2 >>
rect 570300 6400 570900 7400
rect 571900 6400 572500 7400
rect 573500 6400 574100 7400
rect 575100 6400 575700 7400
<< via2 >>
rect 385600 575000 386000 575400
rect 384000 573000 384400 573400
rect 381000 569000 383000 571000
rect 570300 319300 570900 319900
rect 118620 15600 119020 16000
rect 118620 15100 119020 15500
rect 118620 14600 119020 15000
rect 118620 14100 119020 14500
rect 118620 13600 119020 14000
rect 118620 13100 119020 13500
rect 118620 12600 119020 13000
rect 118620 12100 119020 12500
rect 122830 15600 123230 16000
rect 122830 15100 123230 15500
rect 122830 14600 123230 15000
rect 122830 14100 123230 14500
rect 122830 13600 123230 14000
rect 122830 13100 123230 13500
rect 122830 12600 123230 13000
rect 122830 12100 123230 12500
rect 127260 15600 127660 16000
rect 127260 15100 127660 15500
rect 127260 14600 127660 15000
rect 127260 14100 127660 14500
rect 127260 13600 127660 14000
rect 127260 13100 127660 13500
rect 127260 12600 127660 13000
rect 127260 12100 127660 12500
rect 131620 15600 132020 16000
rect 131620 15100 132020 15500
rect 131620 14600 132020 15000
rect 131620 14100 132020 14500
rect 131620 13600 132020 14000
rect 131620 13100 132020 13500
rect 131620 12600 132020 13000
rect 131620 12100 132020 12500
rect 136100 15600 136500 16000
rect 136100 15100 136500 15500
rect 136100 14600 136500 15000
rect 136100 14100 136500 14500
rect 136100 13600 136500 14000
rect 136100 13100 136500 13500
rect 136100 12600 136500 13000
rect 136100 12100 136500 12500
rect 144582 14100 144982 14500
rect 144582 13600 144982 14000
rect 144582 13100 144982 13500
rect 144582 12600 144982 13000
rect 144582 12100 144982 12500
rect 571900 274900 572500 275500
rect 573500 94800 574100 95400
rect 575100 50200 575700 50800
<< metal3 >>
rect 16194 693000 21194 704800
rect 68194 703374 73194 704800
rect 68194 702300 73200 703374
rect 68200 702000 73200 702300
rect 68194 698000 73200 702000
rect 51500 693400 57500 693500
rect 51500 693000 51600 693400
rect 16194 688000 51600 693000
rect 51500 687600 51600 688000
rect 57400 687600 57500 693400
rect 68200 693000 73200 698000
rect 120194 694000 125194 704800
rect 165594 702300 170594 704800
rect 170894 701200 173094 704800
rect 119700 693900 125700 694000
rect 99500 693400 105500 693500
rect 99500 693000 99600 693400
rect 68200 688000 99600 693000
rect 51500 687500 57500 687600
rect 99500 687600 99600 688000
rect 105400 687600 105500 693400
rect 119700 688100 119800 693900
rect 125600 688100 125700 693900
rect 119700 688000 125700 688100
rect 99500 687500 105500 687600
rect 170894 686200 173094 700100
rect 173394 701200 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 173394 698900 175594 700100
rect 222594 701200 224794 704800
rect 173394 698800 179300 698900
rect 173394 696800 177200 698800
rect 179200 696800 179300 698800
rect 173394 696700 179300 696800
rect 222594 686200 224794 700100
rect 225094 701200 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 225094 698900 227294 700100
rect 324294 701200 326494 704800
rect 225094 696700 228700 698900
rect 230900 696700 230910 698900
rect 324294 686200 326494 700100
rect 326794 701200 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 326794 686200 328994 700100
rect 510594 686200 515394 704800
rect 520594 686200 525394 704800
rect 566594 702300 571594 704800
rect 170894 685900 528400 686200
rect 33000 685600 39000 685700
rect 33000 685242 33100 685600
rect -800 680242 33100 685242
rect 33000 679800 33100 680242
rect 38900 685242 39000 685600
rect 38900 680242 39004 685242
rect 170894 681700 524200 685900
rect 528400 681700 528410 685900
rect 536000 682400 540200 682600
rect 536000 681800 536200 682400
rect 536800 681800 537000 682400
rect 537600 681800 537800 682400
rect 538400 681800 538600 682400
rect 539200 681800 539400 682400
rect 540000 682230 540200 682400
rect 582300 682230 584800 682984
rect 540000 681800 584800 682230
rect 170894 681400 528400 681700
rect 536000 681600 584800 681800
rect 536000 681000 536200 681600
rect 536800 681000 537000 681600
rect 537600 681000 537800 681600
rect 538400 681000 538600 681600
rect 539200 681000 539400 681600
rect 540000 681000 584800 681600
rect 536000 680800 584800 681000
rect 38900 679800 39000 680242
rect 33000 679700 39000 679800
rect 536000 680200 536200 680800
rect 536800 680200 537000 680800
rect 537600 680200 537800 680800
rect 538400 680200 538600 680800
rect 539200 680200 539400 680800
rect 540000 680200 584800 680800
rect 536000 680000 584800 680200
rect 536000 679400 536200 680000
rect 536800 679400 537000 680000
rect 537600 679400 537800 680000
rect 538400 679400 538600 680000
rect 539200 679400 539400 680000
rect 540000 679400 584800 680000
rect 536000 679200 584800 679400
rect 536000 678600 536200 679200
rect 536800 678600 537000 679200
rect 537600 678600 537800 679200
rect 538400 678600 538600 679200
rect 539200 678600 539400 679200
rect 540000 678600 584800 679200
rect 536000 678570 584800 678600
rect 536000 678400 540200 678570
rect 582300 677984 584800 678570
rect -800 643842 12000 648642
rect 7200 638642 12000 643842
rect 20000 639600 28000 640000
rect 20000 638642 20400 639600
rect -800 633842 20400 638642
rect 20000 632400 20400 633842
rect 27600 632400 28000 639600
rect 20000 632000 28000 632400
rect 574770 639900 584800 644584
rect 574770 637200 574900 639900
rect 579900 639784 584800 639900
rect 579900 637200 580000 639784
rect 574770 636800 580000 637200
rect 574770 634100 574900 636800
rect 579900 634584 580000 636800
rect 579900 634100 584800 634584
rect 574770 629784 584800 634100
rect 568000 589201 568200 589800
rect 568190 589200 568200 589201
rect 568800 589201 569000 589800
rect 568800 589200 568810 589201
rect 568990 589200 569000 589201
rect 569600 589201 569800 589800
rect 569600 589200 569610 589201
rect 569790 589200 569800 589201
rect 570400 589201 570600 589800
rect 570400 589200 570410 589201
rect 570590 589200 570600 589201
rect 571200 589201 571400 589800
rect 571200 589200 571210 589201
rect 571390 589200 571400 589201
rect 572000 589201 572200 589800
rect 572000 589200 572010 589201
rect 572190 589200 572200 589201
rect 572800 589201 573000 589800
rect 572800 589200 572810 589201
rect 572990 589200 573000 589201
rect 573600 589201 578000 589800
rect 573600 589200 573610 589201
rect 580000 589584 583400 589800
rect 580000 589472 584800 589584
rect 580000 589201 583400 589472
rect 582200 589200 583400 589201
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 544000 583400 544200 584000
rect 544800 583400 545000 584000
rect 545600 583674 583400 584000
rect 545600 583562 584800 583674
rect 545600 583400 583400 583562
rect 385590 575400 386010 575405
rect 385590 575000 385600 575400
rect 386000 575000 555000 575400
rect 555400 575000 555410 575400
rect 385590 574995 386010 575000
rect 383990 573400 384410 573405
rect 383990 573000 384000 573400
rect 384400 573000 553000 573400
rect 553400 573000 553410 573400
rect 383990 572995 384410 573000
rect 380990 571000 383010 571005
rect 380990 569000 381000 571000
rect 383000 569000 550000 571000
rect 552000 569000 552010 571000
rect 380990 568995 383010 569000
rect 7600 567200 12400 567400
rect 7600 564242 7800 567200
rect -800 563800 7800 564242
rect 12200 563800 12400 567200
rect -800 563000 12400 563800
rect -800 559600 7800 563000
rect 12200 559600 12400 563000
rect -800 559442 12400 559600
rect 7600 559400 12400 559442
rect 7664 554242 12336 559400
rect -800 549570 12400 554242
rect 575370 550562 584800 555362
rect -800 549442 1660 549570
rect 575370 545362 580230 550562
rect 497928 540562 584800 545362
rect 469562 533886 477030 534524
rect 900 511870 38001 511890
rect 890 511860 38001 511870
rect 880 511850 38001 511860
rect 870 511840 38001 511850
rect 860 511830 38001 511840
rect 850 511820 38001 511830
rect 840 511810 38001 511820
rect 830 511800 38001 511810
rect 820 511790 38001 511800
rect 810 511780 38001 511790
rect 800 511770 38001 511780
rect 790 511760 38001 511770
rect 780 511750 38001 511760
rect 770 511740 38001 511750
rect 760 511730 38001 511740
rect 750 511720 38001 511730
rect 740 511710 38001 511720
rect 730 511700 38001 511710
rect 720 511690 38001 511700
rect 710 511680 38001 511690
rect 700 511670 38001 511680
rect 690 511660 38001 511670
rect 680 511650 38001 511660
rect 670 511642 38001 511650
rect -800 511530 38001 511642
rect 670 511520 38001 511530
rect 680 511510 38001 511520
rect 690 511500 38001 511510
rect 700 511490 38001 511500
rect 710 511480 38001 511490
rect 720 511470 38001 511480
rect 730 511460 38001 511470
rect 740 511450 38001 511460
rect 750 511440 38001 511450
rect 760 511430 38001 511440
rect 770 511420 38001 511430
rect 780 511410 38001 511420
rect 790 511400 38001 511410
rect 800 511390 38001 511400
rect 810 511380 38001 511390
rect 820 511370 38001 511380
rect 830 511360 38001 511370
rect 840 511350 38001 511360
rect 850 511340 38001 511350
rect 860 511330 38001 511340
rect 870 511320 38001 511330
rect 880 511310 38001 511320
rect 890 511300 38001 511310
rect 900 511290 38001 511300
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect 600 505732 4000 506200
rect -800 505620 4000 505732
rect 600 505200 4000 505620
rect 6000 505200 10000 506200
rect 11000 505200 11200 506200
rect 12200 505200 12400 506200
rect 13400 505200 13600 506200
rect 14600 505200 14800 506200
rect 15800 505200 16000 506200
rect 840 468660 34000 468670
rect 830 468650 34000 468660
rect 820 468640 34000 468650
rect 810 468630 34000 468640
rect 800 468620 34000 468630
rect 790 468610 34000 468620
rect 780 468600 34000 468610
rect 770 468590 34000 468600
rect 760 468580 34000 468590
rect 750 468570 34000 468580
rect 740 468560 34000 468570
rect 730 468550 34000 468560
rect 720 468540 34000 468550
rect 710 468530 34000 468540
rect 700 468520 34000 468530
rect 690 468510 34000 468520
rect 680 468500 34000 468510
rect 670 468490 34000 468500
rect 660 468480 34000 468490
rect 650 468470 34000 468480
rect 640 468460 34000 468470
rect 630 468450 34000 468460
rect 620 468440 34000 468450
rect 610 468430 34000 468440
rect 600 468420 34000 468430
rect -800 468308 34000 468420
rect 600 468300 34000 468308
rect 610 468290 34000 468300
rect 620 468280 34000 468290
rect 630 468270 34000 468280
rect 640 468260 34000 468270
rect 650 468250 34000 468260
rect 660 468240 34000 468250
rect 670 468230 34000 468240
rect 680 468220 34000 468230
rect 690 468210 34000 468220
rect 700 468200 34000 468210
rect 710 468190 34000 468200
rect 720 468180 34000 468190
rect 730 468170 34000 468180
rect 740 468160 34000 468170
rect 750 468150 34000 468160
rect 760 468140 34000 468150
rect 770 468130 34000 468140
rect 780 468120 34000 468130
rect 790 468110 34000 468120
rect 800 468100 34000 468110
rect 810 468090 34000 468100
rect 820 468080 34000 468090
rect 830 468070 34000 468080
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect 600 462510 4000 463000
rect -800 462398 4000 462510
rect 600 462000 4000 462398
rect 6000 462000 10000 463000
rect 11000 462000 11200 463000
rect 12200 462000 12400 463000
rect 13400 462000 13600 463000
rect 14600 462000 14800 463000
rect 15800 462000 16000 463000
rect 840 425440 30000 425450
rect 830 425430 30000 425440
rect 820 425420 30000 425430
rect 810 425410 30000 425420
rect 800 425400 30000 425410
rect 790 425390 30000 425400
rect 780 425380 30000 425390
rect 770 425370 30000 425380
rect 760 425360 30000 425370
rect 750 425350 30000 425360
rect 740 425340 30000 425350
rect 730 425330 30000 425340
rect 720 425320 30000 425330
rect 710 425310 30000 425320
rect 700 425300 30000 425310
rect 690 425290 30000 425300
rect 680 425280 30000 425290
rect 670 425270 30000 425280
rect 660 425260 30000 425270
rect 650 425250 30000 425260
rect 640 425240 30000 425250
rect 630 425230 30000 425240
rect 620 425220 30000 425230
rect 610 425210 30000 425220
rect 600 425198 30000 425210
rect -800 425086 30000 425198
rect 600 425080 30000 425086
rect 610 425070 30000 425080
rect 620 425060 30000 425070
rect 630 425050 30000 425060
rect 640 425040 30000 425050
rect 650 425030 30000 425040
rect 660 425020 30000 425030
rect 670 425010 30000 425020
rect 680 425000 30000 425010
rect 690 424990 30000 425000
rect 700 424980 30000 424990
rect 710 424970 30000 424980
rect 720 424960 30000 424970
rect 730 424950 30000 424960
rect 740 424940 30000 424950
rect 750 424930 30000 424940
rect 760 424920 30000 424930
rect 770 424910 30000 424920
rect 780 424900 30000 424910
rect 790 424890 30000 424900
rect 800 424880 30000 424890
rect 810 424870 30000 424880
rect 820 424860 30000 424870
rect 830 424850 30000 424860
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect 600 419288 4000 419800
rect -800 419176 4000 419288
rect 600 418800 4000 419176
rect 6000 418800 10000 419800
rect 11000 418800 11200 419800
rect 12200 418800 12400 419800
rect 13400 418800 13600 419800
rect 14600 418800 14800 419800
rect 15800 418800 16000 419800
rect 840 382220 26000 382230
rect 830 382210 26000 382220
rect 820 382200 26000 382210
rect 810 382190 26000 382200
rect 800 382180 26000 382190
rect 790 382170 26000 382180
rect 780 382160 26000 382170
rect 770 382150 26000 382160
rect 760 382140 26000 382150
rect 750 382130 26000 382140
rect 740 382120 26000 382130
rect 730 382110 26000 382120
rect 720 382100 26000 382110
rect 710 382090 26000 382100
rect 700 382080 26000 382090
rect 690 382070 26000 382080
rect 680 382060 26000 382070
rect 670 382050 26000 382060
rect 660 382040 26000 382050
rect 650 382030 26000 382040
rect 640 382020 26000 382030
rect 630 382010 26000 382020
rect 620 382000 26000 382010
rect 610 381990 26000 382000
rect 600 381976 26000 381990
rect -800 381864 26000 381976
rect 600 381860 26000 381864
rect 610 381850 26000 381860
rect 620 381840 26000 381850
rect 630 381830 26000 381840
rect 640 381820 26000 381830
rect 650 381810 26000 381820
rect 660 381800 26000 381810
rect 670 381790 26000 381800
rect 680 381780 26000 381790
rect 690 381770 26000 381780
rect 700 381760 26000 381770
rect 710 381750 26000 381760
rect 720 381740 26000 381750
rect 730 381730 26000 381740
rect 740 381720 26000 381730
rect 750 381710 26000 381720
rect 760 381700 26000 381710
rect 770 381690 26000 381700
rect 780 381680 26000 381690
rect 790 381670 26000 381680
rect 800 381660 26000 381670
rect 810 381650 26000 381660
rect 820 381640 26000 381650
rect 830 381630 26000 381640
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect 600 376066 4000 376400
rect -800 375954 4000 376066
rect 600 375400 4000 375954
rect 6000 375400 10000 376400
rect 11000 375400 11200 376400
rect 12200 375400 12400 376400
rect 13400 375400 13600 376400
rect 14600 375400 14800 376400
rect 15800 375400 16000 376400
rect 840 338998 22000 339008
rect 830 338988 22000 338998
rect 820 338978 22000 338988
rect 810 338968 22000 338978
rect 800 338958 22000 338968
rect 790 338948 22000 338958
rect 780 338938 22000 338948
rect 770 338928 22000 338938
rect 760 338918 22000 338928
rect 750 338908 22000 338918
rect 740 338898 22000 338908
rect 730 338888 22000 338898
rect 720 338878 22000 338888
rect 710 338868 22000 338878
rect 700 338858 22000 338868
rect 690 338848 22000 338858
rect 680 338838 22000 338848
rect 670 338828 22000 338838
rect 660 338818 22000 338828
rect 650 338808 22000 338818
rect 640 338798 22000 338808
rect 630 338788 22000 338798
rect 620 338778 22000 338788
rect 610 338768 22000 338778
rect 600 338754 22000 338768
rect -800 338642 22000 338754
rect 600 338638 22000 338642
rect 610 338628 22000 338638
rect 620 338618 22000 338628
rect 630 338608 22000 338618
rect 640 338598 22000 338608
rect 650 338588 22000 338598
rect 660 338578 22000 338588
rect 670 338568 22000 338578
rect 680 338558 22000 338568
rect 690 338548 22000 338558
rect 700 338538 22000 338548
rect 710 338528 22000 338538
rect 720 338518 22000 338528
rect 730 338508 22000 338518
rect 740 338498 22000 338508
rect 750 338488 22000 338498
rect 760 338478 22000 338488
rect 770 338468 22000 338478
rect 780 338458 22000 338468
rect 790 338448 22000 338458
rect 800 338438 22000 338448
rect 810 338428 22000 338438
rect 820 338418 22000 338428
rect 830 338408 22000 338418
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect 600 332844 4000 333200
rect -800 332732 4000 332844
rect 600 332200 4000 332732
rect 6000 332200 10000 333200
rect 11000 332200 11200 333200
rect 12200 332200 12400 333200
rect 13400 332200 13600 333200
rect 14600 332200 14800 333200
rect 15800 332200 16000 333200
rect 20000 331645 22000 338408
rect 24000 335091 26000 381630
rect 28000 339196 30000 424850
rect 32000 342831 34000 468070
rect 36000 452090 38001 511290
rect 469562 486919 470200 533886
rect 471222 528002 476778 528758
rect 536000 528200 540200 528400
rect 536000 528066 536200 528200
rect 471222 488778 471978 528002
rect 526270 527600 536200 528066
rect 536800 527600 537000 528200
rect 537600 527600 537800 528200
rect 538400 527600 538600 528200
rect 539200 527600 539400 528200
rect 540000 527600 540200 528200
rect 526270 527400 540200 527600
rect 526270 526800 536200 527400
rect 536800 526800 537000 527400
rect 537600 526800 537800 527400
rect 538400 526800 538600 527400
rect 539200 526800 539400 527400
rect 540000 526800 540200 527400
rect 526270 526600 540200 526800
rect 526270 526000 536200 526600
rect 536800 526000 537000 526600
rect 537600 526000 537800 526600
rect 538400 526000 538600 526600
rect 539200 526000 539400 526600
rect 540000 526000 540200 526600
rect 526270 525800 540200 526000
rect 526270 525200 536200 525800
rect 536800 525200 537000 525800
rect 537600 525200 537800 525800
rect 538400 525200 538600 525800
rect 539200 525200 539400 525800
rect 540000 525200 540200 525800
rect 526270 525000 540200 525200
rect 526270 524406 536200 525000
rect 536000 524400 536200 524406
rect 536800 524400 537000 525000
rect 537600 524400 537800 525000
rect 538400 524400 538600 525000
rect 539200 524400 539400 525000
rect 540000 524400 540200 525000
rect 536000 524200 540200 524400
rect 473154 522150 477046 523042
rect 473154 490846 474046 522150
rect 474999 516632 477001 517434
rect 474999 493001 475801 516632
rect 544000 514600 545800 514800
rect 544000 514318 544200 514600
rect 530736 514000 544200 514318
rect 544800 514000 545000 514600
rect 545600 514000 545800 514600
rect 530736 513800 546000 514000
rect 530736 513390 544200 513800
rect 544000 513200 544200 513390
rect 544800 513200 545000 513800
rect 545600 513200 546000 513800
rect 544000 513000 546000 513200
rect 481598 494400 482324 506163
rect 497076 505395 498406 507215
rect 524200 505600 528400 505800
rect 524200 505395 524400 505600
rect 497076 505000 524400 505395
rect 525000 505000 525200 505600
rect 525800 505000 526000 505600
rect 526600 505000 526800 505600
rect 527400 505000 527600 505600
rect 528200 505000 528400 505600
rect 497076 504800 528400 505000
rect 497076 504200 524400 504800
rect 525000 504200 525200 504800
rect 525800 504200 526000 504800
rect 526600 504200 526800 504800
rect 527400 504200 527600 504800
rect 528200 504200 528400 504800
rect 497076 504000 528400 504200
rect 497076 503400 524400 504000
rect 525000 503400 525200 504000
rect 525800 503400 526000 504000
rect 526600 503400 526800 504000
rect 527400 503400 527600 504000
rect 528200 503400 528400 504000
rect 497076 503200 528400 503400
rect 497076 502600 524400 503200
rect 525000 502600 525200 503200
rect 525800 502600 526000 503200
rect 526600 502600 526800 503200
rect 527400 502600 527600 503200
rect 528200 502600 528400 503200
rect 497076 502400 528400 502600
rect 497076 502000 524400 502400
rect 524200 501800 524400 502000
rect 525000 501800 525200 502400
rect 525800 501800 526000 502400
rect 526600 501800 526800 502400
rect 527400 501800 527600 502400
rect 528200 501800 528400 502400
rect 524200 501600 528400 501800
rect 568000 499801 568200 500400
rect 568190 499800 568200 499801
rect 568800 499801 569000 500400
rect 568800 499800 568810 499801
rect 568990 499800 569000 499801
rect 569600 499801 569800 500400
rect 569600 499800 569610 499801
rect 569790 499800 569800 499801
rect 570400 499801 570600 500400
rect 570400 499800 570410 499801
rect 570590 499800 570600 499801
rect 571200 499801 571400 500400
rect 571200 499800 571210 499801
rect 571390 499800 571400 499801
rect 572000 499801 572200 500400
rect 572000 499800 572010 499801
rect 572190 499800 572200 499801
rect 572800 499801 573000 500400
rect 572800 499800 572810 499801
rect 572990 499800 573000 499801
rect 573600 499801 578000 500400
rect 573600 499800 573610 499801
rect 580000 500162 583400 500400
rect 580000 500050 584800 500162
rect 580000 499801 583400 500050
rect 582200 499800 583400 499801
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 481598 494252 583400 494400
rect 481598 494140 584800 494252
rect 481598 494001 583400 494140
rect 583000 494000 583400 494001
rect 548000 493001 549000 493100
rect 474999 493000 549000 493001
rect 474999 492200 548100 493000
rect 548900 492200 549000 493000
rect 474999 492199 549000 492200
rect 548000 492100 549000 492199
rect 546000 490846 547000 490900
rect 473154 490800 547000 490846
rect 473154 490000 546100 490800
rect 546900 490000 547000 490800
rect 473154 489954 547000 490000
rect 546000 489900 547000 489954
rect 544000 488800 545000 488900
rect 544000 488778 544100 488800
rect 471222 488022 544100 488778
rect 544000 488000 544100 488022
rect 544900 488000 545000 488800
rect 544000 487900 545000 488000
rect 542000 487000 543000 487100
rect 542000 486919 542100 487000
rect 469562 486281 542100 486919
rect 542000 486200 542100 486281
rect 542900 486200 543000 487000
rect 542000 486100 543000 486200
rect 568000 455401 568200 456000
rect 568190 455400 568200 455401
rect 568800 455401 569000 456000
rect 568800 455400 568810 455401
rect 568990 455400 569000 455401
rect 569600 455401 569800 456000
rect 569600 455400 569610 455401
rect 569790 455400 569800 455401
rect 570400 455401 570600 456000
rect 570400 455400 570410 455401
rect 570590 455400 570600 455401
rect 571200 455401 571400 456000
rect 571200 455400 571210 455401
rect 571390 455400 571400 455401
rect 572000 455401 572200 456000
rect 572000 455400 572010 455401
rect 572190 455400 572200 455401
rect 572800 455401 573000 456000
rect 572800 455400 572810 455401
rect 572990 455400 573000 455401
rect 573600 455401 578000 456000
rect 573600 455400 573610 455401
rect 580000 455740 583400 456000
rect 580000 455628 584800 455740
rect 580000 455401 583400 455628
rect 582200 455400 583400 455401
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 36000 346320 38000 452090
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 554990 449600 555000 450000
rect 555400 449830 583400 450000
rect 555400 449718 584800 449830
rect 555400 449600 583400 449718
rect 568000 411001 568200 411600
rect 568190 411000 568200 411001
rect 568800 411001 569000 411600
rect 568800 411000 568810 411001
rect 568990 411000 569000 411001
rect 569600 411001 569800 411600
rect 569600 411000 569610 411001
rect 569790 411000 569800 411001
rect 570400 411001 570600 411600
rect 570400 411000 570410 411001
rect 570590 411000 570600 411001
rect 571200 411001 571400 411600
rect 571200 411000 571210 411001
rect 571390 411000 571400 411001
rect 572000 411001 572200 411600
rect 572000 411000 572010 411001
rect 572190 411000 572200 411001
rect 572800 411001 573000 411600
rect 572800 411000 572810 411001
rect 572990 411000 573000 411001
rect 573600 411001 578000 411600
rect 573600 411000 573610 411001
rect 580000 411318 583400 411600
rect 580000 411206 584800 411318
rect 580000 411001 583400 411206
rect 582200 411000 583400 411001
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 552990 405200 553000 405600
rect 553400 405408 583400 405600
rect 553400 405296 584800 405408
rect 553400 405200 583400 405296
rect 568000 364601 568200 365200
rect 568190 364600 568200 364601
rect 568800 364601 569000 365200
rect 568800 364600 568810 364601
rect 568990 364600 569000 364601
rect 569600 364601 569800 365200
rect 569600 364600 569610 364601
rect 569790 364600 569800 364601
rect 570400 364601 570600 365200
rect 570400 364600 570410 364601
rect 570590 364600 570600 364601
rect 571200 364601 571400 365200
rect 571200 364600 571210 364601
rect 571390 364600 571400 364601
rect 572000 364601 572200 365200
rect 572000 364600 572010 364601
rect 572190 364600 572200 364601
rect 572800 364601 573000 365200
rect 572800 364600 572810 364601
rect 572990 364600 573000 364601
rect 573600 364601 578000 365200
rect 573600 364600 573610 364601
rect 580000 364896 583400 365200
rect 580000 364784 584800 364896
rect 580000 364601 583400 364784
rect 582200 364600 583400 364601
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 549990 357800 550000 359800
rect 552000 358986 583200 359800
rect 552000 358874 584800 358986
rect 552000 357800 583200 358874
rect 60040 346320 62770 346325
rect 36000 346300 62770 346320
rect 36000 345740 60100 346300
rect 60660 345740 60800 346300
rect 61360 345740 61500 346300
rect 62060 345740 62200 346300
rect 62760 345740 62770 346300
rect 36000 345600 62770 345740
rect 36000 345040 60100 345600
rect 60660 345040 60800 345600
rect 61360 345040 61500 345600
rect 62060 345040 62200 345600
rect 62760 345040 62770 345600
rect 36000 344900 62770 345040
rect 36000 344340 60100 344900
rect 60660 344340 60800 344900
rect 61360 344340 61500 344900
rect 62060 344340 62200 344900
rect 62760 344340 62770 344900
rect 36000 344320 62770 344340
rect 60680 344310 60780 344320
rect 60012 342831 62742 342839
rect 32000 342814 62742 342831
rect 32000 342254 60072 342814
rect 60632 342254 60772 342814
rect 61332 342254 61472 342814
rect 62032 342254 62172 342814
rect 62732 342254 62742 342814
rect 32000 342114 62742 342254
rect 32000 341554 60072 342114
rect 60632 341554 60772 342114
rect 61332 341554 61472 342114
rect 62032 341554 62172 342114
rect 62732 341554 62742 342114
rect 32000 341414 62742 341554
rect 32000 340854 60072 341414
rect 60632 340854 60772 341414
rect 61332 340854 61472 341414
rect 62032 340854 62172 341414
rect 62732 340854 62742 341414
rect 32000 340834 62742 340854
rect 32000 340831 62313 340834
rect 60652 340824 60752 340831
rect 60080 339196 62810 339199
rect 28000 339174 62810 339196
rect 28000 338614 60140 339174
rect 60700 338614 60840 339174
rect 61400 338614 61540 339174
rect 62100 338614 62240 339174
rect 62800 338614 62810 339174
rect 28000 338474 62810 338614
rect 28000 337914 60140 338474
rect 60700 337914 60840 338474
rect 61400 337914 61540 338474
rect 62100 337914 62240 338474
rect 62800 337914 62810 338474
rect 28000 337774 62810 337914
rect 28000 337214 60140 337774
rect 60700 337214 60840 337774
rect 61400 337214 61540 337774
rect 62100 337214 62240 337774
rect 62800 337214 62810 337774
rect 28000 337196 62810 337214
rect 60120 337194 62810 337196
rect 60720 337184 60820 337194
rect 60080 335091 62810 335095
rect 24000 335070 62810 335091
rect 24000 334510 60140 335070
rect 60700 334510 60840 335070
rect 61400 334510 61540 335070
rect 62100 334510 62240 335070
rect 62800 334510 62810 335070
rect 24000 334370 62810 334510
rect 24000 333810 60140 334370
rect 60700 333810 60840 334370
rect 61400 333810 61540 334370
rect 62100 333810 62240 334370
rect 62800 333810 62810 334370
rect 24000 333670 62810 333810
rect 24000 333110 60140 333670
rect 60700 333110 60840 333670
rect 61400 333110 61540 333670
rect 62100 333110 62240 333670
rect 62800 333110 62810 333670
rect 24000 333091 62810 333110
rect 60120 333090 62810 333091
rect 60720 333080 60820 333090
rect 60080 331645 62810 331649
rect 20000 331624 62810 331645
rect 20000 331064 60140 331624
rect 60700 331064 60840 331624
rect 61400 331064 61540 331624
rect 62100 331064 62240 331624
rect 62800 331064 62810 331624
rect 20000 330924 62810 331064
rect 20000 330364 60140 330924
rect 60700 330364 60840 330924
rect 61400 330364 61540 330924
rect 62100 330364 62240 330924
rect 62800 330364 62810 330924
rect 20000 330224 62810 330364
rect 20000 329664 60140 330224
rect 60700 329664 60840 330224
rect 61400 329664 61540 330224
rect 62100 329664 62240 330224
rect 62800 329664 62810 330224
rect 20000 329645 62810 329664
rect 60120 329644 62810 329645
rect 60720 329634 60820 329644
rect 22012 321571 110376 321580
rect 22012 321271 107516 321571
rect 107816 321271 107876 321571
rect 108176 321271 108236 321571
rect 108536 321271 108596 321571
rect 108896 321271 108956 321571
rect 109256 321271 109316 321571
rect 109616 321271 109676 321571
rect 109976 321271 110036 321571
rect 110336 321271 110376 321571
rect 22012 321211 110376 321271
rect 22012 320911 107516 321211
rect 107816 320911 107876 321211
rect 108176 320911 108236 321211
rect 108536 320911 108596 321211
rect 108896 320911 108956 321211
rect 109256 320911 109316 321211
rect 109616 320911 109676 321211
rect 109976 320911 110036 321211
rect 110336 320911 110376 321211
rect 22012 320851 110376 320911
rect 22012 320551 107516 320851
rect 107816 320551 107876 320851
rect 108176 320551 108236 320851
rect 108536 320551 108596 320851
rect 108896 320551 108956 320851
rect 109256 320551 109316 320851
rect 109616 320551 109676 320851
rect 109976 320551 110036 320851
rect 110336 320551 110376 320851
rect 22012 320491 110376 320551
rect 22012 320191 107516 320491
rect 107816 320191 107876 320491
rect 108176 320191 108236 320491
rect 108536 320191 108596 320491
rect 108896 320191 108956 320491
rect 109256 320191 109316 320491
rect 109616 320191 109676 320491
rect 109976 320191 110036 320491
rect 110336 320191 110376 320491
rect 22012 320131 110376 320191
rect 22012 319831 107516 320131
rect 107816 319831 107876 320131
rect 108176 319831 108236 320131
rect 108536 319831 108596 320131
rect 108896 319831 108956 320131
rect 109256 319831 109316 320131
rect 109616 319831 109676 320131
rect 109976 319831 110036 320131
rect 110336 319831 110376 320131
rect 22012 319771 110376 319831
rect 22012 319580 107516 319771
rect 22012 295780 24012 319580
rect 107508 319471 107516 319580
rect 107816 319471 107876 319771
rect 108176 319471 108236 319771
rect 108536 319471 108596 319771
rect 108896 319471 108956 319771
rect 109256 319471 109316 319771
rect 109616 319471 109676 319771
rect 109976 319471 110036 319771
rect 110336 319471 110376 319771
rect 107508 319451 110376 319471
rect 570290 319900 570910 319905
rect 570290 319300 570300 319900
rect 570900 319674 583400 319900
rect 570900 319562 584800 319674
rect 570900 319300 583400 319562
rect 570290 319295 570910 319300
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 840 295770 24012 295780
rect 830 295760 24012 295770
rect 820 295750 24012 295760
rect 810 295740 24012 295750
rect 800 295730 24012 295740
rect 790 295720 24012 295730
rect 780 295710 24012 295720
rect 770 295700 24012 295710
rect 760 295690 24012 295700
rect 750 295680 24012 295690
rect 740 295670 24012 295680
rect 730 295660 24012 295670
rect 720 295650 24012 295660
rect 710 295640 24012 295650
rect 700 295630 24012 295640
rect 690 295620 24012 295630
rect 680 295610 24012 295620
rect 670 295600 24012 295610
rect 660 295590 24012 295600
rect 650 295580 24012 295590
rect 640 295570 24012 295580
rect 630 295560 24012 295570
rect 620 295550 24012 295560
rect 610 295540 24012 295550
rect 600 295532 24012 295540
rect -800 295420 24012 295532
rect 600 295410 24012 295420
rect 610 295400 24012 295410
rect 620 295390 24012 295400
rect 630 295380 24012 295390
rect 640 295370 24012 295380
rect 650 295360 24012 295370
rect 660 295350 24012 295360
rect 670 295340 24012 295350
rect 680 295330 24012 295340
rect 690 295320 24012 295330
rect 700 295310 24012 295320
rect 710 295300 24012 295310
rect 720 295290 24012 295300
rect 730 295280 24012 295290
rect 740 295270 24012 295280
rect 750 295260 24012 295270
rect 760 295250 24012 295260
rect 770 295240 24012 295250
rect 780 295230 24012 295240
rect 790 295220 24012 295230
rect 800 295210 24012 295220
rect 810 295200 24012 295210
rect 820 295190 24012 295200
rect 830 295180 24012 295190
rect 26012 315880 188772 315889
rect 26012 315580 185912 315880
rect 186212 315580 186272 315880
rect 186572 315580 186632 315880
rect 186932 315580 186992 315880
rect 187292 315580 187352 315880
rect 187652 315580 187712 315880
rect 188012 315580 188072 315880
rect 188372 315580 188432 315880
rect 188732 315580 188772 315880
rect 547990 315600 548000 316600
rect 549000 316128 583400 316600
rect 549000 316016 584800 316128
rect 549000 315600 583400 316016
rect 26012 315520 188772 315580
rect 26012 315220 185912 315520
rect 186212 315220 186272 315520
rect 186572 315220 186632 315520
rect 186932 315220 186992 315520
rect 187292 315220 187352 315520
rect 187652 315220 187712 315520
rect 188012 315220 188072 315520
rect 188372 315220 188432 315520
rect 188732 315220 188772 315520
rect 26012 315160 188772 315220
rect 26012 314860 185912 315160
rect 186212 314860 186272 315160
rect 186572 314860 186632 315160
rect 186932 314860 186992 315160
rect 187292 314860 187352 315160
rect 187652 314860 187712 315160
rect 188012 314860 188072 315160
rect 188372 314860 188432 315160
rect 188732 314860 188772 315160
rect 26012 314800 188772 314860
rect 583520 314834 584800 314946
rect 26012 314500 185912 314800
rect 186212 314500 186272 314800
rect 186572 314500 186632 314800
rect 186932 314500 186992 314800
rect 187292 314500 187352 314800
rect 187652 314500 187712 314800
rect 188012 314500 188072 314800
rect 188372 314500 188432 314800
rect 188732 314500 188772 314800
rect 26012 314440 188772 314500
rect 26012 314140 185912 314440
rect 186212 314140 186272 314440
rect 186572 314140 186632 314440
rect 186932 314140 186992 314440
rect 187292 314140 187352 314440
rect 187652 314140 187712 314440
rect 188012 314140 188072 314440
rect 188372 314140 188432 314440
rect 188732 314140 188772 314440
rect 26012 314080 188772 314140
rect 26012 313889 185912 314080
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect 600 289622 4000 290000
rect -800 289510 4000 289622
rect 600 289000 4000 289510
rect 6000 289000 10000 290000
rect 11000 289000 11200 290000
rect 12200 289000 12400 290000
rect 13400 289000 13600 290000
rect 14600 289000 14800 290000
rect 15800 289000 16000 290000
rect 26012 252760 28012 313889
rect 185892 313780 185912 313889
rect 186212 313780 186272 314080
rect 186572 313780 186632 314080
rect 186932 313780 186992 314080
rect 187292 313780 187352 314080
rect 187652 313780 187712 314080
rect 188012 313780 188072 314080
rect 188372 313780 188432 314080
rect 188732 313780 188772 314080
rect 185892 313760 188772 313780
rect 583520 313652 584800 313764
rect 840 252750 28012 252760
rect 830 252740 28012 252750
rect 820 252730 28012 252740
rect 810 252720 28012 252730
rect 800 252710 28012 252720
rect 790 252700 28012 252710
rect 780 252690 28012 252700
rect 770 252680 28012 252690
rect 760 252670 28012 252680
rect 750 252660 28012 252670
rect 740 252650 28012 252660
rect 730 252640 28012 252650
rect 720 252630 28012 252640
rect 710 252620 28012 252630
rect 700 252610 28012 252620
rect 690 252600 28012 252610
rect 680 252590 28012 252600
rect 670 252580 28012 252590
rect 660 252570 28012 252580
rect 650 252560 28012 252570
rect 640 252550 28012 252560
rect 630 252540 28012 252550
rect 620 252530 28012 252540
rect 610 252520 28012 252530
rect 600 252510 28012 252520
rect -800 252398 28012 252510
rect 600 252390 28012 252398
rect 610 252380 28012 252390
rect 620 252370 28012 252380
rect 630 252360 28012 252370
rect 640 252350 28012 252360
rect 650 252340 28012 252350
rect 660 252330 28012 252340
rect 670 252320 28012 252330
rect 680 252310 28012 252320
rect 690 252300 28012 252310
rect 700 252290 28012 252300
rect 710 252280 28012 252290
rect 720 252270 28012 252280
rect 730 252260 28012 252270
rect 740 252250 28012 252260
rect 750 252240 28012 252250
rect 760 252230 28012 252240
rect 770 252220 28012 252230
rect 780 252210 28012 252220
rect 790 252200 28012 252210
rect 800 252190 28012 252200
rect 810 252180 28012 252190
rect 820 252170 28012 252180
rect 830 252160 28012 252170
rect 30012 310414 264594 310423
rect 30012 310114 261734 310414
rect 262034 310114 262094 310414
rect 262394 310114 262454 310414
rect 262754 310114 262814 310414
rect 263114 310114 263174 310414
rect 263474 310114 263534 310414
rect 263834 310114 263894 310414
rect 264194 310114 264254 310414
rect 264554 310114 264594 310414
rect 30012 310054 264594 310114
rect 30012 309754 261734 310054
rect 262034 309754 262094 310054
rect 262394 309754 262454 310054
rect 262754 309754 262814 310054
rect 263114 309754 263174 310054
rect 263474 309754 263534 310054
rect 263834 309754 263894 310054
rect 264194 309754 264254 310054
rect 264554 309754 264594 310054
rect 30012 309694 264594 309754
rect 30012 309394 261734 309694
rect 262034 309394 262094 309694
rect 262394 309394 262454 309694
rect 262754 309394 262814 309694
rect 263114 309394 263174 309694
rect 263474 309394 263534 309694
rect 263834 309394 263894 309694
rect 264194 309394 264254 309694
rect 264554 309394 264594 309694
rect 30012 309334 264594 309394
rect 30012 309034 261734 309334
rect 262034 309034 262094 309334
rect 262394 309034 262454 309334
rect 262754 309034 262814 309334
rect 263114 309034 263174 309334
rect 263474 309034 263534 309334
rect 263834 309034 263894 309334
rect 264194 309034 264254 309334
rect 264554 309034 264594 309334
rect 30012 308974 264594 309034
rect 30012 308674 261734 308974
rect 262034 308674 262094 308974
rect 262394 308674 262454 308974
rect 262754 308674 262814 308974
rect 263114 308674 263174 308974
rect 263474 308674 263534 308974
rect 263834 308674 263894 308974
rect 264194 308674 264254 308974
rect 264554 308674 264594 308974
rect 30012 308614 264594 308674
rect 30012 308423 261734 308614
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect 600 246600 4000 247000
rect -800 246488 4000 246600
rect 600 246000 4000 246488
rect 6000 246000 10000 247000
rect 11000 246000 11200 247000
rect 12200 246000 12400 247000
rect 13400 246000 13600 247000
rect 14600 246000 14800 247000
rect 15800 246000 16000 247000
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 3000 178800 11000 179200
rect 3000 177688 3400 178800
rect -800 172888 3400 177688
rect 3000 171600 3400 172888
rect 10600 171600 11000 178800
rect 3000 171200 11000 171600
rect 4600 167688 9400 171200
rect -800 162888 9400 167688
rect 30012 125140 32012 308423
rect 261726 308314 261734 308423
rect 262034 308314 262094 308614
rect 262394 308314 262454 308614
rect 262754 308314 262814 308614
rect 263114 308314 263174 308614
rect 263474 308314 263534 308614
rect 263834 308314 263894 308614
rect 264194 308314 264254 308614
rect 264554 308314 264594 308614
rect 261726 308294 264594 308314
rect 840 125130 32012 125140
rect 830 125120 32012 125130
rect 820 125110 32012 125120
rect 810 125100 32012 125110
rect 800 125090 32012 125100
rect 790 125080 32012 125090
rect 780 125070 32012 125080
rect 770 125060 32012 125070
rect 760 125050 32012 125060
rect 750 125040 32012 125050
rect 740 125030 32012 125040
rect 730 125020 32012 125030
rect 720 125010 32012 125020
rect 710 125000 32012 125010
rect 700 124990 32012 125000
rect 690 124980 32012 124990
rect 680 124970 32012 124980
rect 670 124960 32012 124970
rect 660 124950 32012 124960
rect 650 124940 32012 124950
rect 640 124930 32012 124940
rect 630 124920 32012 124930
rect 620 124910 32012 124920
rect 610 124900 32012 124910
rect 600 124888 32012 124900
rect -800 124776 32012 124888
rect 600 124770 32012 124776
rect 610 124760 32012 124770
rect 620 124750 32012 124760
rect 630 124740 32012 124750
rect 640 124730 32012 124740
rect 650 124720 32012 124730
rect 660 124710 32012 124720
rect 670 124700 32012 124710
rect 680 124690 32012 124700
rect 690 124680 32012 124690
rect 700 124670 32012 124680
rect 710 124660 32012 124670
rect 720 124650 32012 124660
rect 730 124640 32012 124650
rect 740 124630 32012 124640
rect 750 124620 32012 124630
rect 760 124610 32012 124620
rect 770 124600 32012 124610
rect 780 124590 32012 124600
rect 790 124580 32012 124590
rect 800 124570 32012 124580
rect 810 124560 32012 124570
rect 820 124550 32012 124560
rect 830 124540 32012 124550
rect 34012 304188 342392 304197
rect 34012 303888 339528 304188
rect 339828 303888 339888 304188
rect 340188 303888 340248 304188
rect 340548 303888 340608 304188
rect 340908 303888 340968 304188
rect 341268 303888 341328 304188
rect 341628 303888 341688 304188
rect 341988 303888 342048 304188
rect 342348 303888 342392 304188
rect 34012 303828 342392 303888
rect 34012 303528 339528 303828
rect 339828 303528 339888 303828
rect 340188 303528 340248 303828
rect 340548 303528 340608 303828
rect 340908 303528 340968 303828
rect 341268 303528 341328 303828
rect 341628 303528 341688 303828
rect 341988 303528 342048 303828
rect 342348 303528 342392 303828
rect 34012 303468 342392 303528
rect 34012 303168 339528 303468
rect 339828 303168 339888 303468
rect 340188 303168 340248 303468
rect 340548 303168 340608 303468
rect 340908 303168 340968 303468
rect 341268 303168 341328 303468
rect 341628 303168 341688 303468
rect 341988 303168 342048 303468
rect 342348 303168 342392 303468
rect 34012 303108 342392 303168
rect 34012 302808 339528 303108
rect 339828 302808 339888 303108
rect 340188 302808 340248 303108
rect 340548 302808 340608 303108
rect 340908 302808 340968 303108
rect 341268 302808 341328 303108
rect 341628 302808 341688 303108
rect 341988 302808 342048 303108
rect 342348 302808 342392 303108
rect 34012 302748 342392 302808
rect 34012 302448 339528 302748
rect 339828 302448 339888 302748
rect 340188 302448 340248 302748
rect 340548 302448 340608 302748
rect 340908 302448 340968 302748
rect 341268 302448 341328 302748
rect 341628 302448 341688 302748
rect 341988 302448 342048 302748
rect 342348 302448 342392 302748
rect 34012 302388 342392 302448
rect 34012 302197 339528 302388
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect 600 118978 4000 119400
rect -800 118866 4000 118978
rect 600 118400 4000 118866
rect 6000 118400 10000 119400
rect 11000 118400 11200 119400
rect 12200 118400 12400 119400
rect 13400 118400 13600 119400
rect 14600 118400 14800 119400
rect 15800 118400 16000 119400
rect 34012 81920 36012 302197
rect 339520 302088 339528 302197
rect 339828 302088 339888 302388
rect 340188 302088 340248 302388
rect 340548 302088 340608 302388
rect 340908 302088 340968 302388
rect 341268 302088 341328 302388
rect 341628 302088 341688 302388
rect 341988 302088 342048 302388
rect 342348 302197 342392 302388
rect 342348 302088 342388 302197
rect 339520 302068 342388 302088
rect 571890 275500 572510 275505
rect 571890 274900 571900 275500
rect 572500 275252 583400 275500
rect 572500 275140 584800 275252
rect 572500 274900 583400 275140
rect 571890 274895 572510 274900
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 545990 271200 546000 272200
rect 547000 271706 583400 272200
rect 547000 271594 584800 271706
rect 547000 271200 583400 271594
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect 573490 95400 574110 95405
rect 573490 94800 573500 95400
rect 574100 95230 583400 95400
rect 574100 95118 584800 95230
rect 574100 94800 583400 95118
rect 573490 94795 574110 94800
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 543990 91200 544000 92200
rect 545000 91684 583200 92200
rect 545000 91572 584800 91684
rect 545000 91200 583200 91572
rect 840 81910 36012 81920
rect 830 81900 36012 81910
rect 820 81890 36012 81900
rect 810 81880 36012 81890
rect 800 81870 36012 81880
rect 790 81860 36012 81870
rect 780 81850 36012 81860
rect 770 81840 36012 81850
rect 760 81830 36012 81840
rect 750 81820 36012 81830
rect 740 81810 36012 81820
rect 730 81800 36012 81810
rect 720 81790 36012 81800
rect 710 81780 36012 81790
rect 700 81770 36012 81780
rect 690 81760 36012 81770
rect 680 81750 36012 81760
rect 670 81740 36012 81750
rect 660 81730 36012 81740
rect 650 81720 36012 81730
rect 640 81710 36012 81720
rect 630 81700 36012 81710
rect 620 81690 36012 81700
rect 610 81680 36012 81690
rect 600 81666 36012 81680
rect -800 81554 36012 81666
rect 600 81550 36012 81554
rect 610 81540 36012 81550
rect 620 81530 36012 81540
rect 630 81520 36012 81530
rect 640 81510 36012 81520
rect 650 81500 36012 81510
rect 660 81490 36012 81500
rect 670 81480 36012 81490
rect 680 81470 36012 81480
rect 690 81460 36012 81470
rect 700 81450 36012 81460
rect 710 81440 36012 81450
rect 720 81430 36012 81440
rect 730 81420 36012 81430
rect 740 81410 36012 81420
rect 750 81400 36012 81410
rect 760 81390 36012 81400
rect 770 81380 36012 81390
rect 780 81370 36012 81380
rect 790 81360 36012 81370
rect 800 81350 36012 81360
rect 810 81340 36012 81350
rect 820 81330 36012 81340
rect 830 81320 36012 81330
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect 600 75756 4000 76200
rect -800 75644 4000 75756
rect 600 75200 4000 75644
rect 6000 75200 10000 76200
rect 11000 75200 11200 76200
rect 12200 75200 12400 76200
rect 13400 75200 13600 76200
rect 14600 75200 14800 76200
rect 15800 75200 16000 76200
rect 575090 50800 575710 50805
rect 575090 50200 575100 50800
rect 575700 50572 583400 50800
rect 575700 50460 584800 50572
rect 575700 50200 583400 50460
rect 575090 50195 575710 50200
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 541990 46400 542000 47400
rect 543000 47026 583400 47400
rect 543000 46914 584800 47026
rect 543000 46400 583400 46914
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect 840 35140 139200 35150
rect 830 35130 139200 35140
rect 820 35120 139200 35130
rect 810 35110 139200 35120
rect 800 35100 139200 35110
rect 790 35090 139200 35100
rect 780 35080 139200 35090
rect 770 35070 139200 35080
rect 760 35060 139200 35070
rect 750 35050 139200 35060
rect 740 35040 139200 35050
rect 730 35030 139200 35040
rect 720 35020 139200 35030
rect 710 35010 139200 35020
rect 700 35000 139200 35010
rect 690 34990 139200 35000
rect 680 34980 139200 34990
rect 670 34970 139200 34980
rect 660 34960 139200 34970
rect 650 34950 139200 34960
rect 640 34940 139200 34950
rect 630 34930 139200 34940
rect 620 34920 139200 34930
rect 610 34910 139200 34920
rect 600 34898 139200 34910
rect -800 34786 139200 34898
rect 600 34780 139200 34786
rect 610 34770 139200 34780
rect 620 34760 139200 34770
rect 630 34750 139200 34760
rect 640 34740 139200 34750
rect 650 34730 139200 34740
rect 660 34720 139200 34730
rect 670 34710 139200 34720
rect 680 34700 139200 34710
rect 690 34690 139200 34700
rect 700 34680 139200 34690
rect 710 34670 139200 34680
rect 720 34660 139200 34670
rect 730 34650 139200 34660
rect 740 34640 139200 34650
rect 750 34630 139200 34640
rect 760 34620 139200 34630
rect 770 34610 139200 34620
rect 780 34600 139200 34610
rect 790 34590 139200 34600
rect 800 34580 139200 34590
rect 810 34570 139200 34580
rect 820 34560 139200 34570
rect 830 34550 139200 34560
rect 139800 34550 139960 35150
rect 140560 34550 140740 35150
rect 141340 34550 141500 35150
rect 142100 34550 142155 35150
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 118590 15580 118600 16020
rect 119040 15580 119050 16020
rect 122800 15580 122810 16020
rect 123250 15580 123260 16020
rect 127230 15580 127240 16020
rect 127680 15580 127690 16020
rect 131590 15580 131600 16020
rect 132040 15580 132050 16020
rect 136070 15580 136080 16020
rect 136520 15580 136530 16020
rect 583520 15728 584800 15840
rect 118590 15080 118600 15520
rect 119040 15080 119050 15520
rect 122800 15080 122810 15520
rect 123250 15080 123260 15520
rect 127230 15080 127240 15520
rect 127680 15080 127690 15520
rect 131590 15080 131600 15520
rect 132040 15080 132050 15520
rect 136070 15080 136080 15520
rect 136520 15080 136530 15520
rect -800 14546 480 14658
rect 118590 14580 118600 15020
rect 119040 14580 119050 15020
rect 122800 14580 122810 15020
rect 123250 14580 123260 15020
rect 127230 14580 127240 15020
rect 127680 14580 127690 15020
rect 131590 14580 131600 15020
rect 132040 14580 132050 15020
rect 136070 14580 136080 15020
rect 136520 14580 136530 15020
rect 583520 14546 584800 14658
rect 118590 14080 118600 14520
rect 119040 14080 119050 14520
rect 122800 14080 122810 14520
rect 123250 14080 123260 14520
rect 127230 14080 127240 14520
rect 127680 14080 127690 14520
rect 131590 14080 131600 14520
rect 132040 14080 132050 14520
rect 136070 14080 136080 14520
rect 136520 14080 136530 14520
rect 144552 14080 144562 14520
rect 145002 14080 145012 14520
rect 118590 13580 118600 14020
rect 119040 13580 119050 14020
rect 122800 13580 122810 14020
rect 123250 13580 123260 14020
rect 127230 13580 127240 14020
rect 127680 13580 127690 14020
rect 131590 13580 131600 14020
rect 132040 13580 132050 14020
rect 136070 13580 136080 14020
rect 136520 13580 136530 14020
rect 144552 13580 144562 14020
rect 145002 13580 145012 14020
rect -800 13364 480 13476
rect 118590 13080 118600 13520
rect 119040 13080 119050 13520
rect 122800 13080 122810 13520
rect 123250 13080 123260 13520
rect 127230 13080 127240 13520
rect 127680 13080 127690 13520
rect 131590 13080 131600 13520
rect 132040 13080 132050 13520
rect 136070 13080 136080 13520
rect 136520 13080 136530 13520
rect 144552 13080 144562 13520
rect 145002 13080 145012 13520
rect 583520 13364 584800 13476
rect 118590 12580 118600 13020
rect 119040 12580 119050 13020
rect 122800 12580 122810 13020
rect 123250 12580 123260 13020
rect 127230 12580 127240 13020
rect 127680 12580 127690 13020
rect 131590 12580 131600 13020
rect 132040 12580 132050 13020
rect 136070 12580 136080 13020
rect 136520 12580 136530 13020
rect 144552 12580 144562 13020
rect 145002 12580 145012 13020
rect -800 12182 480 12294
rect 118590 12080 118600 12520
rect 119040 12080 119050 12520
rect 122800 12080 122810 12520
rect 123250 12080 123260 12520
rect 127230 12080 127240 12520
rect 127680 12080 127690 12520
rect 131590 12080 131600 12520
rect 132040 12080 132050 12520
rect 136070 12080 136080 12520
rect 136520 12080 136530 12520
rect 144552 12080 144562 12520
rect 145002 12080 145012 12520
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 170894 700100 173094 701200
rect 173394 700100 175594 701200
rect 222594 700100 224794 701200
rect 225094 700100 227294 701200
rect 324294 700100 326494 701200
rect 326794 700100 328994 701200
rect 578000 589200 580000 589800
rect 4000 505200 6000 506200
rect 4000 462000 6000 463000
rect 4000 418800 6000 419800
rect 4000 375400 6000 376400
rect 4000 332200 6000 333200
rect 578000 499800 580000 500400
rect 578000 455400 580000 456000
rect 578000 411000 580000 411600
rect 578000 364600 580000 365200
rect 4000 289000 6000 290000
rect 4000 246000 6000 247000
rect 4000 118400 6000 119400
rect 4000 75200 6000 76200
<< via3 >>
rect 51600 687600 57400 693400
rect 99600 687600 105400 693400
rect 119800 688100 125600 693900
rect 177200 696800 179200 698800
rect 228700 696700 230900 698900
rect 33100 679800 38900 685600
rect 524200 681700 528400 685900
rect 536200 681800 536800 682400
rect 537000 681800 537600 682400
rect 537800 681800 538400 682400
rect 538600 681800 539200 682400
rect 539400 681800 540000 682400
rect 536200 681000 536800 681600
rect 537000 681000 537600 681600
rect 537800 681000 538400 681600
rect 538600 681000 539200 681600
rect 539400 681000 540000 681600
rect 536200 680200 536800 680800
rect 537000 680200 537600 680800
rect 537800 680200 538400 680800
rect 538600 680200 539200 680800
rect 539400 680200 540000 680800
rect 536200 679400 536800 680000
rect 537000 679400 537600 680000
rect 537800 679400 538400 680000
rect 538600 679400 539200 680000
rect 539400 679400 540000 680000
rect 536200 678600 536800 679200
rect 537000 678600 537600 679200
rect 537800 678600 538400 679200
rect 538600 678600 539200 679200
rect 539400 678600 540000 679200
rect 20400 632400 27600 639600
rect 574900 637200 579900 639900
rect 574900 634100 579900 636800
rect 568200 589200 568800 589800
rect 569000 589200 569600 589800
rect 569800 589200 570400 589800
rect 570600 589200 571200 589800
rect 571400 589200 572000 589800
rect 572200 589200 572800 589800
rect 573000 589200 573600 589800
rect 544200 583400 544800 584000
rect 545000 583400 545600 584000
rect 555000 575000 555400 575400
rect 553000 573000 553400 573400
rect 550000 569000 552000 571000
rect 7800 563800 12200 567200
rect 7800 559600 12200 563000
rect 10000 505200 11000 506200
rect 11200 505200 12200 506200
rect 12400 505200 13400 506200
rect 13600 505200 14600 506200
rect 14800 505200 15800 506200
rect 10000 462000 11000 463000
rect 11200 462000 12200 463000
rect 12400 462000 13400 463000
rect 13600 462000 14600 463000
rect 14800 462000 15800 463000
rect 10000 418800 11000 419800
rect 11200 418800 12200 419800
rect 12400 418800 13400 419800
rect 13600 418800 14600 419800
rect 14800 418800 15800 419800
rect 10000 375400 11000 376400
rect 11200 375400 12200 376400
rect 12400 375400 13400 376400
rect 13600 375400 14600 376400
rect 14800 375400 15800 376400
rect 10000 332200 11000 333200
rect 11200 332200 12200 333200
rect 12400 332200 13400 333200
rect 13600 332200 14600 333200
rect 14800 332200 15800 333200
rect 536200 527600 536800 528200
rect 537000 527600 537600 528200
rect 537800 527600 538400 528200
rect 538600 527600 539200 528200
rect 539400 527600 540000 528200
rect 536200 526800 536800 527400
rect 537000 526800 537600 527400
rect 537800 526800 538400 527400
rect 538600 526800 539200 527400
rect 539400 526800 540000 527400
rect 536200 526000 536800 526600
rect 537000 526000 537600 526600
rect 537800 526000 538400 526600
rect 538600 526000 539200 526600
rect 539400 526000 540000 526600
rect 536200 525200 536800 525800
rect 537000 525200 537600 525800
rect 537800 525200 538400 525800
rect 538600 525200 539200 525800
rect 539400 525200 540000 525800
rect 536200 524400 536800 525000
rect 537000 524400 537600 525000
rect 537800 524400 538400 525000
rect 538600 524400 539200 525000
rect 539400 524400 540000 525000
rect 544200 514000 544800 514600
rect 545000 514000 545600 514600
rect 544200 513200 544800 513800
rect 545000 513200 545600 513800
rect 524400 505000 525000 505600
rect 525200 505000 525800 505600
rect 526000 505000 526600 505600
rect 526800 505000 527400 505600
rect 527600 505000 528200 505600
rect 524400 504200 525000 504800
rect 525200 504200 525800 504800
rect 526000 504200 526600 504800
rect 526800 504200 527400 504800
rect 527600 504200 528200 504800
rect 524400 503400 525000 504000
rect 525200 503400 525800 504000
rect 526000 503400 526600 504000
rect 526800 503400 527400 504000
rect 527600 503400 528200 504000
rect 524400 502600 525000 503200
rect 525200 502600 525800 503200
rect 526000 502600 526600 503200
rect 526800 502600 527400 503200
rect 527600 502600 528200 503200
rect 524400 501800 525000 502400
rect 525200 501800 525800 502400
rect 526000 501800 526600 502400
rect 526800 501800 527400 502400
rect 527600 501800 528200 502400
rect 568200 499800 568800 500400
rect 569000 499800 569600 500400
rect 569800 499800 570400 500400
rect 570600 499800 571200 500400
rect 571400 499800 572000 500400
rect 572200 499800 572800 500400
rect 573000 499800 573600 500400
rect 548100 492200 548900 493000
rect 546100 490000 546900 490800
rect 544100 488000 544900 488800
rect 542100 486200 542900 487000
rect 568200 455400 568800 456000
rect 569000 455400 569600 456000
rect 569800 455400 570400 456000
rect 570600 455400 571200 456000
rect 571400 455400 572000 456000
rect 572200 455400 572800 456000
rect 573000 455400 573600 456000
rect 555000 449600 555400 450000
rect 568200 411000 568800 411600
rect 569000 411000 569600 411600
rect 569800 411000 570400 411600
rect 570600 411000 571200 411600
rect 571400 411000 572000 411600
rect 572200 411000 572800 411600
rect 573000 411000 573600 411600
rect 553000 405200 553400 405600
rect 568200 364600 568800 365200
rect 569000 364600 569600 365200
rect 569800 364600 570400 365200
rect 570600 364600 571200 365200
rect 571400 364600 572000 365200
rect 572200 364600 572800 365200
rect 573000 364600 573600 365200
rect 550000 357800 552000 359800
rect 60100 345740 60660 346300
rect 60800 345740 61360 346300
rect 61500 345740 62060 346300
rect 62200 345740 62760 346300
rect 60100 345040 60660 345600
rect 60800 345040 61360 345600
rect 61500 345040 62060 345600
rect 62200 345040 62760 345600
rect 60100 344340 60660 344900
rect 60800 344340 61360 344900
rect 61500 344340 62060 344900
rect 62200 344340 62760 344900
rect 60072 342254 60632 342814
rect 60772 342254 61332 342814
rect 61472 342254 62032 342814
rect 62172 342254 62732 342814
rect 60072 341554 60632 342114
rect 60772 341554 61332 342114
rect 61472 341554 62032 342114
rect 62172 341554 62732 342114
rect 60072 340854 60632 341414
rect 60772 340854 61332 341414
rect 61472 340854 62032 341414
rect 62172 340854 62732 341414
rect 60140 338614 60700 339174
rect 60840 338614 61400 339174
rect 61540 338614 62100 339174
rect 62240 338614 62800 339174
rect 60140 337914 60700 338474
rect 60840 337914 61400 338474
rect 61540 337914 62100 338474
rect 62240 337914 62800 338474
rect 60140 337214 60700 337774
rect 60840 337214 61400 337774
rect 61540 337214 62100 337774
rect 62240 337214 62800 337774
rect 60140 334510 60700 335070
rect 60840 334510 61400 335070
rect 61540 334510 62100 335070
rect 62240 334510 62800 335070
rect 60140 333810 60700 334370
rect 60840 333810 61400 334370
rect 61540 333810 62100 334370
rect 62240 333810 62800 334370
rect 60140 333110 60700 333670
rect 60840 333110 61400 333670
rect 61540 333110 62100 333670
rect 62240 333110 62800 333670
rect 60140 331064 60700 331624
rect 60840 331064 61400 331624
rect 61540 331064 62100 331624
rect 62240 331064 62800 331624
rect 60140 330364 60700 330924
rect 60840 330364 61400 330924
rect 61540 330364 62100 330924
rect 62240 330364 62800 330924
rect 60140 329664 60700 330224
rect 60840 329664 61400 330224
rect 61540 329664 62100 330224
rect 62240 329664 62800 330224
rect 107516 321271 107816 321571
rect 107876 321271 108176 321571
rect 108236 321271 108536 321571
rect 108596 321271 108896 321571
rect 108956 321271 109256 321571
rect 109316 321271 109616 321571
rect 109676 321271 109976 321571
rect 110036 321271 110336 321571
rect 107516 320911 107816 321211
rect 107876 320911 108176 321211
rect 108236 320911 108536 321211
rect 108596 320911 108896 321211
rect 108956 320911 109256 321211
rect 109316 320911 109616 321211
rect 109676 320911 109976 321211
rect 110036 320911 110336 321211
rect 107516 320551 107816 320851
rect 107876 320551 108176 320851
rect 108236 320551 108536 320851
rect 108596 320551 108896 320851
rect 108956 320551 109256 320851
rect 109316 320551 109616 320851
rect 109676 320551 109976 320851
rect 110036 320551 110336 320851
rect 107516 320191 107816 320491
rect 107876 320191 108176 320491
rect 108236 320191 108536 320491
rect 108596 320191 108896 320491
rect 108956 320191 109256 320491
rect 109316 320191 109616 320491
rect 109676 320191 109976 320491
rect 110036 320191 110336 320491
rect 107516 319831 107816 320131
rect 107876 319831 108176 320131
rect 108236 319831 108536 320131
rect 108596 319831 108896 320131
rect 108956 319831 109256 320131
rect 109316 319831 109616 320131
rect 109676 319831 109976 320131
rect 110036 319831 110336 320131
rect 107516 319471 107816 319771
rect 107876 319471 108176 319771
rect 108236 319471 108536 319771
rect 108596 319471 108896 319771
rect 108956 319471 109256 319771
rect 109316 319471 109616 319771
rect 109676 319471 109976 319771
rect 110036 319471 110336 319771
rect 185912 315580 186212 315880
rect 186272 315580 186572 315880
rect 186632 315580 186932 315880
rect 186992 315580 187292 315880
rect 187352 315580 187652 315880
rect 187712 315580 188012 315880
rect 188072 315580 188372 315880
rect 188432 315580 188732 315880
rect 548000 315600 549000 316600
rect 185912 315220 186212 315520
rect 186272 315220 186572 315520
rect 186632 315220 186932 315520
rect 186992 315220 187292 315520
rect 187352 315220 187652 315520
rect 187712 315220 188012 315520
rect 188072 315220 188372 315520
rect 188432 315220 188732 315520
rect 185912 314860 186212 315160
rect 186272 314860 186572 315160
rect 186632 314860 186932 315160
rect 186992 314860 187292 315160
rect 187352 314860 187652 315160
rect 187712 314860 188012 315160
rect 188072 314860 188372 315160
rect 188432 314860 188732 315160
rect 185912 314500 186212 314800
rect 186272 314500 186572 314800
rect 186632 314500 186932 314800
rect 186992 314500 187292 314800
rect 187352 314500 187652 314800
rect 187712 314500 188012 314800
rect 188072 314500 188372 314800
rect 188432 314500 188732 314800
rect 185912 314140 186212 314440
rect 186272 314140 186572 314440
rect 186632 314140 186932 314440
rect 186992 314140 187292 314440
rect 187352 314140 187652 314440
rect 187712 314140 188012 314440
rect 188072 314140 188372 314440
rect 188432 314140 188732 314440
rect 10000 289000 11000 290000
rect 11200 289000 12200 290000
rect 12400 289000 13400 290000
rect 13600 289000 14600 290000
rect 14800 289000 15800 290000
rect 185912 313780 186212 314080
rect 186272 313780 186572 314080
rect 186632 313780 186932 314080
rect 186992 313780 187292 314080
rect 187352 313780 187652 314080
rect 187712 313780 188012 314080
rect 188072 313780 188372 314080
rect 188432 313780 188732 314080
rect 261734 310114 262034 310414
rect 262094 310114 262394 310414
rect 262454 310114 262754 310414
rect 262814 310114 263114 310414
rect 263174 310114 263474 310414
rect 263534 310114 263834 310414
rect 263894 310114 264194 310414
rect 264254 310114 264554 310414
rect 261734 309754 262034 310054
rect 262094 309754 262394 310054
rect 262454 309754 262754 310054
rect 262814 309754 263114 310054
rect 263174 309754 263474 310054
rect 263534 309754 263834 310054
rect 263894 309754 264194 310054
rect 264254 309754 264554 310054
rect 261734 309394 262034 309694
rect 262094 309394 262394 309694
rect 262454 309394 262754 309694
rect 262814 309394 263114 309694
rect 263174 309394 263474 309694
rect 263534 309394 263834 309694
rect 263894 309394 264194 309694
rect 264254 309394 264554 309694
rect 261734 309034 262034 309334
rect 262094 309034 262394 309334
rect 262454 309034 262754 309334
rect 262814 309034 263114 309334
rect 263174 309034 263474 309334
rect 263534 309034 263834 309334
rect 263894 309034 264194 309334
rect 264254 309034 264554 309334
rect 261734 308674 262034 308974
rect 262094 308674 262394 308974
rect 262454 308674 262754 308974
rect 262814 308674 263114 308974
rect 263174 308674 263474 308974
rect 263534 308674 263834 308974
rect 263894 308674 264194 308974
rect 264254 308674 264554 308974
rect 10000 246000 11000 247000
rect 11200 246000 12200 247000
rect 12400 246000 13400 247000
rect 13600 246000 14600 247000
rect 14800 246000 15800 247000
rect 3400 171600 10600 178800
rect 261734 308314 262034 308614
rect 262094 308314 262394 308614
rect 262454 308314 262754 308614
rect 262814 308314 263114 308614
rect 263174 308314 263474 308614
rect 263534 308314 263834 308614
rect 263894 308314 264194 308614
rect 264254 308314 264554 308614
rect 339528 303888 339828 304188
rect 339888 303888 340188 304188
rect 340248 303888 340548 304188
rect 340608 303888 340908 304188
rect 340968 303888 341268 304188
rect 341328 303888 341628 304188
rect 341688 303888 341988 304188
rect 342048 303888 342348 304188
rect 339528 303528 339828 303828
rect 339888 303528 340188 303828
rect 340248 303528 340548 303828
rect 340608 303528 340908 303828
rect 340968 303528 341268 303828
rect 341328 303528 341628 303828
rect 341688 303528 341988 303828
rect 342048 303528 342348 303828
rect 339528 303168 339828 303468
rect 339888 303168 340188 303468
rect 340248 303168 340548 303468
rect 340608 303168 340908 303468
rect 340968 303168 341268 303468
rect 341328 303168 341628 303468
rect 341688 303168 341988 303468
rect 342048 303168 342348 303468
rect 339528 302808 339828 303108
rect 339888 302808 340188 303108
rect 340248 302808 340548 303108
rect 340608 302808 340908 303108
rect 340968 302808 341268 303108
rect 341328 302808 341628 303108
rect 341688 302808 341988 303108
rect 342048 302808 342348 303108
rect 339528 302448 339828 302748
rect 339888 302448 340188 302748
rect 340248 302448 340548 302748
rect 340608 302448 340908 302748
rect 340968 302448 341268 302748
rect 341328 302448 341628 302748
rect 341688 302448 341988 302748
rect 342048 302448 342348 302748
rect 10000 118400 11000 119400
rect 11200 118400 12200 119400
rect 12400 118400 13400 119400
rect 13600 118400 14600 119400
rect 14800 118400 15800 119400
rect 339528 302088 339828 302388
rect 339888 302088 340188 302388
rect 340248 302088 340548 302388
rect 340608 302088 340908 302388
rect 340968 302088 341268 302388
rect 341328 302088 341628 302388
rect 341688 302088 341988 302388
rect 342048 302088 342348 302388
rect 546000 271200 547000 272200
rect 544000 91200 545000 92200
rect 10000 75200 11000 76200
rect 11200 75200 12200 76200
rect 12400 75200 13400 76200
rect 13600 75200 14600 76200
rect 14800 75200 15800 76200
rect 542000 46400 543000 47400
rect 139200 34550 139800 35150
rect 139960 34550 140560 35150
rect 140740 34550 141340 35150
rect 141500 34550 142100 35150
rect 118600 16000 119040 16020
rect 118600 15600 118620 16000
rect 118620 15600 119020 16000
rect 119020 15600 119040 16000
rect 118600 15580 119040 15600
rect 122810 16000 123250 16020
rect 122810 15600 122830 16000
rect 122830 15600 123230 16000
rect 123230 15600 123250 16000
rect 122810 15580 123250 15600
rect 127240 16000 127680 16020
rect 127240 15600 127260 16000
rect 127260 15600 127660 16000
rect 127660 15600 127680 16000
rect 127240 15580 127680 15600
rect 131600 16000 132040 16020
rect 131600 15600 131620 16000
rect 131620 15600 132020 16000
rect 132020 15600 132040 16000
rect 131600 15580 132040 15600
rect 136080 16000 136520 16020
rect 136080 15600 136100 16000
rect 136100 15600 136500 16000
rect 136500 15600 136520 16000
rect 136080 15580 136520 15600
rect 118600 15500 119040 15520
rect 118600 15100 118620 15500
rect 118620 15100 119020 15500
rect 119020 15100 119040 15500
rect 118600 15080 119040 15100
rect 122810 15500 123250 15520
rect 122810 15100 122830 15500
rect 122830 15100 123230 15500
rect 123230 15100 123250 15500
rect 122810 15080 123250 15100
rect 127240 15500 127680 15520
rect 127240 15100 127260 15500
rect 127260 15100 127660 15500
rect 127660 15100 127680 15500
rect 127240 15080 127680 15100
rect 131600 15500 132040 15520
rect 131600 15100 131620 15500
rect 131620 15100 132020 15500
rect 132020 15100 132040 15500
rect 131600 15080 132040 15100
rect 136080 15500 136520 15520
rect 136080 15100 136100 15500
rect 136100 15100 136500 15500
rect 136500 15100 136520 15500
rect 136080 15080 136520 15100
rect 118600 15000 119040 15020
rect 118600 14600 118620 15000
rect 118620 14600 119020 15000
rect 119020 14600 119040 15000
rect 118600 14580 119040 14600
rect 122810 15000 123250 15020
rect 122810 14600 122830 15000
rect 122830 14600 123230 15000
rect 123230 14600 123250 15000
rect 122810 14580 123250 14600
rect 127240 15000 127680 15020
rect 127240 14600 127260 15000
rect 127260 14600 127660 15000
rect 127660 14600 127680 15000
rect 127240 14580 127680 14600
rect 131600 15000 132040 15020
rect 131600 14600 131620 15000
rect 131620 14600 132020 15000
rect 132020 14600 132040 15000
rect 131600 14580 132040 14600
rect 136080 15000 136520 15020
rect 136080 14600 136100 15000
rect 136100 14600 136500 15000
rect 136500 14600 136520 15000
rect 136080 14580 136520 14600
rect 118600 14500 119040 14520
rect 118600 14100 118620 14500
rect 118620 14100 119020 14500
rect 119020 14100 119040 14500
rect 118600 14080 119040 14100
rect 122810 14500 123250 14520
rect 122810 14100 122830 14500
rect 122830 14100 123230 14500
rect 123230 14100 123250 14500
rect 122810 14080 123250 14100
rect 127240 14500 127680 14520
rect 127240 14100 127260 14500
rect 127260 14100 127660 14500
rect 127660 14100 127680 14500
rect 127240 14080 127680 14100
rect 131600 14500 132040 14520
rect 131600 14100 131620 14500
rect 131620 14100 132020 14500
rect 132020 14100 132040 14500
rect 131600 14080 132040 14100
rect 136080 14500 136520 14520
rect 136080 14100 136100 14500
rect 136100 14100 136500 14500
rect 136500 14100 136520 14500
rect 136080 14080 136520 14100
rect 144562 14500 145002 14520
rect 144562 14100 144582 14500
rect 144582 14100 144982 14500
rect 144982 14100 145002 14500
rect 144562 14080 145002 14100
rect 118600 14000 119040 14020
rect 118600 13600 118620 14000
rect 118620 13600 119020 14000
rect 119020 13600 119040 14000
rect 118600 13580 119040 13600
rect 122810 14000 123250 14020
rect 122810 13600 122830 14000
rect 122830 13600 123230 14000
rect 123230 13600 123250 14000
rect 122810 13580 123250 13600
rect 127240 14000 127680 14020
rect 127240 13600 127260 14000
rect 127260 13600 127660 14000
rect 127660 13600 127680 14000
rect 127240 13580 127680 13600
rect 131600 14000 132040 14020
rect 131600 13600 131620 14000
rect 131620 13600 132020 14000
rect 132020 13600 132040 14000
rect 131600 13580 132040 13600
rect 136080 14000 136520 14020
rect 136080 13600 136100 14000
rect 136100 13600 136500 14000
rect 136500 13600 136520 14000
rect 136080 13580 136520 13600
rect 144562 14000 145002 14020
rect 144562 13600 144582 14000
rect 144582 13600 144982 14000
rect 144982 13600 145002 14000
rect 144562 13580 145002 13600
rect 118600 13500 119040 13520
rect 118600 13100 118620 13500
rect 118620 13100 119020 13500
rect 119020 13100 119040 13500
rect 118600 13080 119040 13100
rect 122810 13500 123250 13520
rect 122810 13100 122830 13500
rect 122830 13100 123230 13500
rect 123230 13100 123250 13500
rect 122810 13080 123250 13100
rect 127240 13500 127680 13520
rect 127240 13100 127260 13500
rect 127260 13100 127660 13500
rect 127660 13100 127680 13500
rect 127240 13080 127680 13100
rect 131600 13500 132040 13520
rect 131600 13100 131620 13500
rect 131620 13100 132020 13500
rect 132020 13100 132040 13500
rect 131600 13080 132040 13100
rect 136080 13500 136520 13520
rect 136080 13100 136100 13500
rect 136100 13100 136500 13500
rect 136500 13100 136520 13500
rect 136080 13080 136520 13100
rect 144562 13500 145002 13520
rect 144562 13100 144582 13500
rect 144582 13100 144982 13500
rect 144982 13100 145002 13500
rect 144562 13080 145002 13100
rect 118600 13000 119040 13020
rect 118600 12600 118620 13000
rect 118620 12600 119020 13000
rect 119020 12600 119040 13000
rect 118600 12580 119040 12600
rect 122810 13000 123250 13020
rect 122810 12600 122830 13000
rect 122830 12600 123230 13000
rect 123230 12600 123250 13000
rect 122810 12580 123250 12600
rect 127240 13000 127680 13020
rect 127240 12600 127260 13000
rect 127260 12600 127660 13000
rect 127660 12600 127680 13000
rect 127240 12580 127680 12600
rect 131600 13000 132040 13020
rect 131600 12600 131620 13000
rect 131620 12600 132020 13000
rect 132020 12600 132040 13000
rect 131600 12580 132040 12600
rect 136080 13000 136520 13020
rect 136080 12600 136100 13000
rect 136100 12600 136500 13000
rect 136500 12600 136520 13000
rect 136080 12580 136520 12600
rect 144562 13000 145002 13020
rect 144562 12600 144582 13000
rect 144582 12600 144982 13000
rect 144982 12600 145002 13000
rect 144562 12580 145002 12600
rect 118600 12500 119040 12520
rect 118600 12100 118620 12500
rect 118620 12100 119020 12500
rect 119020 12100 119040 12500
rect 118600 12080 119040 12100
rect 122810 12500 123250 12520
rect 122810 12100 122830 12500
rect 122830 12100 123230 12500
rect 123230 12100 123250 12500
rect 122810 12080 123250 12100
rect 127240 12500 127680 12520
rect 127240 12100 127260 12500
rect 127260 12100 127660 12500
rect 127660 12100 127680 12500
rect 127240 12080 127680 12100
rect 131600 12500 132040 12520
rect 131600 12100 131620 12500
rect 131620 12100 132020 12500
rect 132020 12100 132040 12500
rect 131600 12080 132040 12100
rect 136080 12500 136520 12520
rect 136080 12100 136100 12500
rect 136100 12100 136500 12500
rect 136500 12100 136520 12500
rect 136080 12080 136520 12100
rect 144562 12500 145002 12520
rect 144562 12100 144582 12500
rect 144582 12100 144982 12500
rect 144982 12100 145002 12500
rect 144562 12080 145002 12100
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 119700 693900 125700 694000
rect 51500 693400 57500 693500
rect 51500 687600 51600 693400
rect 57400 687600 57500 693400
rect 51500 687500 57500 687600
rect 99500 693400 105500 693500
rect 99500 687600 99600 693400
rect 105400 687600 105500 693400
rect 119700 688100 119800 693900
rect 125600 688100 125700 693900
rect 119700 688000 125700 688100
rect 99500 687500 105500 687600
rect 33000 685600 39000 685700
rect 33000 679800 33100 685600
rect 38900 679800 39000 685600
rect 33000 679700 39000 679800
rect 20000 639600 28000 640000
rect 20000 632400 20400 639600
rect 27600 632400 28000 639600
rect 20000 632000 28000 632400
rect 21000 529000 27000 632000
rect 34000 538000 38000 679700
rect 52000 548500 57000 687500
rect 100000 560500 105000 687500
rect 120194 572500 125194 688000
rect 524200 685901 528400 686200
rect 524199 685900 528401 685901
rect 524199 681700 524200 685900
rect 528400 681700 528401 685900
rect 524199 681699 528401 681700
rect 536000 682400 540200 682600
rect 536000 681800 536200 682400
rect 536800 681800 537000 682400
rect 537600 681800 537800 682400
rect 538400 681800 538600 682400
rect 539200 681800 539400 682400
rect 540000 681800 540200 682400
rect 524200 679300 528400 681699
rect 120194 567500 299500 572500
rect 100000 555500 221700 560500
rect 52000 543500 145900 548500
rect 34000 534000 67000 538000
rect 140900 533500 145900 543500
rect 216700 535500 221700 555500
rect 294500 533500 299500 567500
rect 389500 567200 397500 606640
rect 389500 560200 389600 567200
rect 397400 559600 397500 567200
rect 389600 559400 397500 559600
rect 20000 528800 28000 529000
rect 20000 521200 20200 528800
rect 27800 521200 28000 528800
rect 20000 521000 28000 521200
rect 34000 511800 42000 512000
rect 9999 506200 11001 506201
rect 9999 505200 10000 506200
rect 11000 505200 11001 506200
rect 9999 505199 11001 505200
rect 11199 506200 12201 506201
rect 11199 505200 11200 506200
rect 12200 505200 12201 506200
rect 11199 505199 12201 505200
rect 12399 506200 13401 506201
rect 12399 505200 12400 506200
rect 13400 505200 13401 506200
rect 12399 505199 13401 505200
rect 13599 506200 14601 506201
rect 13599 505200 13600 506200
rect 14600 505200 14601 506200
rect 13599 505199 14601 505200
rect 14799 506200 15801 506201
rect 14799 505200 14800 506200
rect 15800 505200 15801 506200
rect 14799 505199 15801 505200
rect 34000 504200 34200 511800
rect 41800 504200 42000 511800
rect 524200 505800 528400 677300
rect 536000 681600 540200 681800
rect 536000 681000 536200 681600
rect 536800 681000 537000 681600
rect 537600 681000 537800 681600
rect 538400 681000 538600 681600
rect 539200 681000 539400 681600
rect 540000 681000 540200 681600
rect 536000 680800 540200 681000
rect 536000 680200 536200 680800
rect 536800 680200 537000 680800
rect 537600 680200 537800 680800
rect 538400 680200 538600 680800
rect 539200 680200 539400 680800
rect 540000 680200 540200 680800
rect 536000 680000 540200 680200
rect 536000 679400 536200 680000
rect 536800 679400 537000 680000
rect 537600 679400 537800 680000
rect 538400 679400 538600 680000
rect 539200 679400 539400 680000
rect 540000 679400 540200 680000
rect 536000 679200 540200 679400
rect 536000 678600 536200 679200
rect 536800 678600 537000 679200
rect 537600 678600 537800 679200
rect 538400 678600 538600 679200
rect 539200 678600 539400 679200
rect 540000 678600 540200 679200
rect 536000 528200 540200 678600
rect 568000 639900 580000 640000
rect 568000 637200 574900 639900
rect 579900 637200 580000 639900
rect 568000 636800 580000 637200
rect 568000 634100 574900 636800
rect 579900 634100 580000 636800
rect 568000 634000 580000 634100
rect 568000 589800 574000 634000
rect 568000 589200 568200 589800
rect 568800 589200 569000 589800
rect 569600 589200 569800 589800
rect 570400 589200 570600 589800
rect 571200 589200 571400 589800
rect 572000 589200 572200 589800
rect 572800 589200 573000 589800
rect 573600 589200 574000 589800
rect 536000 527600 536200 528200
rect 536800 527600 537000 528200
rect 537600 527600 537800 528200
rect 538400 527600 538600 528200
rect 539200 527600 539400 528200
rect 540000 527600 540200 528200
rect 536000 527400 540200 527600
rect 536000 526800 536200 527400
rect 536800 526800 537000 527400
rect 537600 526800 537800 527400
rect 538400 526800 538600 527400
rect 539200 526800 539400 527400
rect 540000 526800 540200 527400
rect 536000 526600 540200 526800
rect 536000 526000 536200 526600
rect 536800 526000 537000 526600
rect 537600 526000 537800 526600
rect 538400 526000 538600 526600
rect 539200 526000 539400 526600
rect 540000 526000 540200 526600
rect 536000 525800 540200 526000
rect 536000 525200 536200 525800
rect 536800 525200 537000 525800
rect 537600 525200 537800 525800
rect 538400 525200 538600 525800
rect 539200 525200 539400 525800
rect 540000 525200 540200 525800
rect 536000 525000 540200 525200
rect 536000 524400 536200 525000
rect 536800 524400 537000 525000
rect 537600 524400 537800 525000
rect 538400 524400 538600 525000
rect 539200 524400 539400 525000
rect 540000 524400 540200 525000
rect 536000 524200 540200 524400
rect 544000 584000 546000 584200
rect 544000 583400 544200 584000
rect 544800 583400 545000 584000
rect 545600 583400 546000 584000
rect 544000 514600 546000 583400
rect 554999 575400 555401 575401
rect 554999 575000 555000 575400
rect 555400 575000 555401 575400
rect 554999 574999 555401 575000
rect 552999 573400 553401 573401
rect 552999 573000 553000 573400
rect 553400 573000 553401 573400
rect 552999 572999 553401 573000
rect 549999 571000 552001 571001
rect 549999 569000 550000 571000
rect 552000 569000 552001 571000
rect 549999 568999 552001 569000
rect 544000 514000 544200 514600
rect 544800 514000 545000 514600
rect 545600 514000 546000 514600
rect 544000 513800 546000 514000
rect 544000 513200 544200 513800
rect 544800 513200 545000 513800
rect 545600 513200 546000 513800
rect 544000 513000 546000 513200
rect 34000 504000 42000 504200
rect 524202 505600 528398 505800
rect 524202 505000 524400 505600
rect 525000 505000 525200 505600
rect 525800 505000 526000 505600
rect 526600 505000 526800 505600
rect 527400 505000 527600 505600
rect 528200 505000 528398 505600
rect 524202 504800 528398 505000
rect 524202 504200 524400 504800
rect 525000 504200 525200 504800
rect 525800 504200 526000 504800
rect 526600 504200 526800 504800
rect 527400 504200 527600 504800
rect 528200 504200 528398 504800
rect 524202 504000 528398 504200
rect 9999 463000 11001 463001
rect 9999 462000 10000 463000
rect 11000 462000 11001 463000
rect 9999 461999 11001 462000
rect 11199 463000 12201 463001
rect 11199 462000 11200 463000
rect 12200 462000 12201 463000
rect 11199 461999 12201 462000
rect 12399 463000 13401 463001
rect 12399 462000 12400 463000
rect 13400 462000 13401 463000
rect 12399 461999 13401 462000
rect 13599 463000 14601 463001
rect 13599 462000 13600 463000
rect 14600 462000 14601 463000
rect 13599 461999 14601 462000
rect 14799 463000 15801 463001
rect 14799 462000 14800 463000
rect 15800 462000 15801 463000
rect 14799 461999 15801 462000
rect 9999 419800 11001 419801
rect 9999 418800 10000 419800
rect 11000 418800 11001 419800
rect 9999 418799 11001 418800
rect 11199 419800 12201 419801
rect 11199 418800 11200 419800
rect 12200 418800 12201 419800
rect 11199 418799 12201 418800
rect 12399 419800 13401 419801
rect 12399 418800 12400 419800
rect 13400 418800 13401 419800
rect 12399 418799 13401 418800
rect 13599 419800 14601 419801
rect 13599 418800 13600 419800
rect 14600 418800 14601 419800
rect 13599 418799 14601 418800
rect 14799 419800 15801 419801
rect 14799 418800 14800 419800
rect 15800 418800 15801 419800
rect 14799 418799 15801 418800
rect 9999 376400 11001 376401
rect 9999 375400 10000 376400
rect 11000 375400 11001 376400
rect 9999 375399 11001 375400
rect 11199 376400 12201 376401
rect 11199 375400 11200 376400
rect 12200 375400 12201 376400
rect 11199 375399 12201 375400
rect 12399 376400 13401 376401
rect 12399 375400 12400 376400
rect 13400 375400 13401 376400
rect 12399 375399 13401 375400
rect 13599 376400 14601 376401
rect 13599 375400 13600 376400
rect 14600 375400 14601 376400
rect 13599 375399 14601 375400
rect 14799 376400 15801 376401
rect 14799 375400 14800 376400
rect 15800 375400 15801 376400
rect 14799 375399 15801 375400
rect 9999 333200 11001 333201
rect 9999 332200 10000 333200
rect 11000 332200 11001 333200
rect 9999 332199 11001 332200
rect 11199 333200 12201 333201
rect 11199 332200 11200 333200
rect 12200 332200 12201 333200
rect 11199 332199 12201 332200
rect 12399 333200 13401 333201
rect 12399 332200 12400 333200
rect 13400 332200 13401 333200
rect 12399 332199 13401 332200
rect 13599 333200 14601 333201
rect 13599 332200 13600 333200
rect 14600 332200 14601 333200
rect 13599 332199 14601 332200
rect 14799 333200 15801 333201
rect 14799 332200 14800 333200
rect 15800 332200 15801 333200
rect 14799 332199 15801 332200
rect 9999 290000 11001 290001
rect 9999 289000 10000 290000
rect 11000 289000 11001 290000
rect 9999 288999 11001 289000
rect 11199 290000 12201 290001
rect 11199 289000 11200 290000
rect 12200 289000 12201 290000
rect 11199 288999 12201 289000
rect 12399 290000 13401 290001
rect 12399 289000 12400 290000
rect 13400 289000 13401 290000
rect 12399 288999 13401 289000
rect 13599 290000 14601 290001
rect 13599 289000 13600 290000
rect 14600 289000 14601 290000
rect 13599 288999 14601 289000
rect 14799 290000 15801 290001
rect 14799 289000 14800 290000
rect 15800 289000 15801 290000
rect 14799 288999 15801 289000
rect 9999 247000 11001 247001
rect 9999 246000 10000 247000
rect 11000 246000 11001 247000
rect 9999 245999 11001 246000
rect 11199 247000 12201 247001
rect 11199 246000 11200 247000
rect 12200 246000 12201 247000
rect 11199 245999 12201 246000
rect 12399 247000 13401 247001
rect 12399 246000 12400 247000
rect 13400 246000 13401 247000
rect 12399 245999 13401 246000
rect 13599 247000 14601 247001
rect 13599 246000 13600 247000
rect 14600 246000 14601 247000
rect 13599 245999 14601 246000
rect 14799 247000 15801 247001
rect 14799 246000 14800 247000
rect 15800 246000 15801 247000
rect 14799 245999 15801 246000
rect 35000 197114 41000 504000
rect 524202 503400 524400 504000
rect 525000 503400 525200 504000
rect 525800 503400 526000 504000
rect 526600 503400 526800 504000
rect 527400 503400 527600 504000
rect 528200 503400 528398 504000
rect 524202 503200 528398 503400
rect 524202 502600 524400 503200
rect 525000 502600 525200 503200
rect 525800 502600 526000 503200
rect 526600 502600 526800 503200
rect 527400 502600 527600 503200
rect 528200 502600 528398 503200
rect 524202 502400 528398 502600
rect 524202 501800 524400 502400
rect 525000 501800 525200 502400
rect 525800 501800 526000 502400
rect 526600 501800 526800 502400
rect 527400 501800 527600 502400
rect 528200 501800 528398 502400
rect 524200 501600 528400 501800
rect 548000 493000 549000 493100
rect 548000 492200 548100 493000
rect 548900 492200 549000 493000
rect 546000 490800 547000 490900
rect 546000 490000 546100 490800
rect 546900 490000 547000 490800
rect 544000 488800 545000 488900
rect 544000 488000 544100 488800
rect 544900 488000 545000 488800
rect 542000 487000 543000 487100
rect 542000 486200 542100 487000
rect 542900 486200 543000 487000
rect 117388 370900 120268 371034
rect 117388 369100 117500 370900
rect 120100 369100 120268 370900
rect 60040 346310 62820 346350
rect 60040 345710 60080 346310
rect 60680 345710 60780 346310
rect 61380 345710 61480 346310
rect 62080 345710 62180 346310
rect 62780 345710 62820 346310
rect 60040 345610 62820 345710
rect 60040 345010 60080 345610
rect 60680 345010 60780 345610
rect 61380 345010 61480 345610
rect 62080 345010 62180 345610
rect 62780 345010 62820 345610
rect 60040 344910 62820 345010
rect 60040 344310 60080 344910
rect 60680 344310 60780 344910
rect 61380 344310 61480 344910
rect 62080 344310 62180 344910
rect 62780 344310 62820 344910
rect 60040 344280 62820 344310
rect 60012 342824 62792 342864
rect 60012 342224 60052 342824
rect 60652 342224 60752 342824
rect 61352 342224 61452 342824
rect 62052 342224 62152 342824
rect 62752 342224 62792 342824
rect 60012 342124 62792 342224
rect 60012 341524 60052 342124
rect 60652 341524 60752 342124
rect 61352 341524 61452 342124
rect 62052 341524 62152 342124
rect 62752 341524 62792 342124
rect 60012 341424 62792 341524
rect 60012 340824 60052 341424
rect 60652 340824 60752 341424
rect 61352 340824 61452 341424
rect 62052 340824 62152 341424
rect 62752 340824 62792 341424
rect 60012 340794 62792 340824
rect 60080 339184 62860 339224
rect 60080 338584 60120 339184
rect 60720 338584 60820 339184
rect 61420 338584 61520 339184
rect 62120 338584 62220 339184
rect 62820 338584 62860 339184
rect 60080 338484 62860 338584
rect 60080 337884 60120 338484
rect 60720 337884 60820 338484
rect 61420 337884 61520 338484
rect 62120 337884 62220 338484
rect 62820 337884 62860 338484
rect 60080 337784 62860 337884
rect 60080 337184 60120 337784
rect 60720 337184 60820 337784
rect 61420 337184 61520 337784
rect 62120 337184 62220 337784
rect 62820 337184 62860 337784
rect 60080 337154 62860 337184
rect 60080 335080 62860 335120
rect 60080 334480 60120 335080
rect 60720 334480 60820 335080
rect 61420 334480 61520 335080
rect 62120 334480 62220 335080
rect 62820 334480 62860 335080
rect 60080 334380 62860 334480
rect 60080 333780 60120 334380
rect 60720 333780 60820 334380
rect 61420 333780 61520 334380
rect 62120 333780 62220 334380
rect 62820 333780 62860 334380
rect 60080 333680 62860 333780
rect 60080 333080 60120 333680
rect 60720 333080 60820 333680
rect 61420 333080 61520 333680
rect 62120 333080 62220 333680
rect 62820 333080 62860 333680
rect 60080 333050 62860 333080
rect 60080 331634 62860 331674
rect 60080 331034 60120 331634
rect 60720 331034 60820 331634
rect 61420 331034 61520 331634
rect 62120 331034 62220 331634
rect 62820 331034 62860 331634
rect 60080 330934 62860 331034
rect 60080 330334 60120 330934
rect 60720 330334 60820 330934
rect 61420 330334 61520 330934
rect 62120 330334 62220 330934
rect 62820 330334 62860 330934
rect 60080 330234 62860 330334
rect 60080 329634 60120 330234
rect 60720 329634 60820 330234
rect 61420 329634 61520 330234
rect 62120 329634 62220 330234
rect 62820 329634 62860 330234
rect 60080 329604 62860 329634
rect 107508 321571 110366 329740
rect 107508 321271 107516 321571
rect 107816 321271 107876 321571
rect 108176 321271 108236 321571
rect 108536 321271 108596 321571
rect 108896 321271 108956 321571
rect 109256 321271 109316 321571
rect 109616 321271 109676 321571
rect 109976 321271 110036 321571
rect 110336 321271 110366 321571
rect 107508 321211 110366 321271
rect 107508 320911 107516 321211
rect 107816 320911 107876 321211
rect 108176 320911 108236 321211
rect 108536 320911 108596 321211
rect 108896 320911 108956 321211
rect 109256 320911 109316 321211
rect 109616 320911 109676 321211
rect 109976 320911 110036 321211
rect 110336 320911 110366 321211
rect 107508 320851 110366 320911
rect 107508 320551 107516 320851
rect 107816 320551 107876 320851
rect 108176 320551 108236 320851
rect 108536 320551 108596 320851
rect 108896 320551 108956 320851
rect 109256 320551 109316 320851
rect 109616 320551 109676 320851
rect 109976 320551 110036 320851
rect 110336 320551 110366 320851
rect 107508 320491 110366 320551
rect 107508 320191 107516 320491
rect 107816 320191 107876 320491
rect 108176 320191 108236 320491
rect 108536 320191 108596 320491
rect 108896 320191 108956 320491
rect 109256 320191 109316 320491
rect 109616 320191 109676 320491
rect 109976 320191 110036 320491
rect 110336 320191 110366 320491
rect 107508 320131 110366 320191
rect 107508 319831 107516 320131
rect 107816 319831 107876 320131
rect 108176 319831 108236 320131
rect 108536 319831 108596 320131
rect 108896 319831 108956 320131
rect 109256 319831 109316 320131
rect 109616 319831 109676 320131
rect 109976 319831 110036 320131
rect 110336 319831 110366 320131
rect 107508 319771 110366 319831
rect 107508 319471 107516 319771
rect 107816 319471 107876 319771
rect 108176 319471 108236 319771
rect 108536 319471 108596 319771
rect 108896 319471 108956 319771
rect 109256 319471 109316 319771
rect 109616 319471 109676 319771
rect 109976 319471 110036 319771
rect 110336 319471 110366 319771
rect 107508 319440 110366 319471
rect 3000 178800 11000 179200
rect 3000 171600 3400 178800
rect 10600 178200 11000 178800
rect 35000 178200 41000 181000
rect 10600 172200 41000 178200
rect 10600 171600 11000 172200
rect 3000 171200 11000 171600
rect 9999 119400 11001 119401
rect 9999 118400 10000 119400
rect 11000 118400 11001 119400
rect 9999 118399 11001 118400
rect 11199 119400 12201 119401
rect 11199 118400 11200 119400
rect 12200 118400 12201 119400
rect 11199 118399 12201 118400
rect 12399 119400 13401 119401
rect 12399 118400 12400 119400
rect 13400 118400 13401 119400
rect 12399 118399 13401 118400
rect 13599 119400 14601 119401
rect 13599 118400 13600 119400
rect 14600 118400 14601 119400
rect 13599 118399 14601 118400
rect 14799 119400 15801 119401
rect 14799 118400 14800 119400
rect 15800 118400 15801 119400
rect 14799 118399 15801 118400
rect 9999 76200 11001 76201
rect 9999 75200 10000 76200
rect 11000 75200 11001 76200
rect 9999 75199 11001 75200
rect 11199 76200 12201 76201
rect 11199 75200 11200 76200
rect 12200 75200 12201 76200
rect 11199 75199 12201 75200
rect 12399 76200 13401 76201
rect 12399 75200 12400 76200
rect 13400 75200 13401 76200
rect 12399 75199 13401 75200
rect 13599 76200 14601 76201
rect 13599 75200 13600 76200
rect 14600 75200 14601 76200
rect 13599 75199 14601 75200
rect 14799 76200 15801 76201
rect 14799 75200 14800 76200
rect 15800 75200 15801 76200
rect 14799 75199 15801 75200
rect 117388 16020 120268 369100
rect 142709 334351 145430 369926
rect 117388 15580 118600 16020
rect 119040 15580 120268 16020
rect 117388 15520 120268 15580
rect 117388 15080 118600 15520
rect 119040 15080 120268 15520
rect 117388 15020 120268 15080
rect 117388 14580 118600 15020
rect 119040 14580 120268 15020
rect 117388 14520 120268 14580
rect 117388 14080 118600 14520
rect 119040 14080 120268 14520
rect 117388 14020 120268 14080
rect 117388 13580 118600 14020
rect 119040 13580 120268 14020
rect 117388 13520 120268 13580
rect 117388 13080 118600 13520
rect 119040 13080 120268 13520
rect 117388 13020 120268 13080
rect 117388 12580 118600 13020
rect 119040 12580 120268 13020
rect 117388 12520 120268 12580
rect 117388 12080 118600 12520
rect 119040 12080 120268 12520
rect 117388 12000 120268 12080
rect 121706 331726 145430 334351
rect 121706 331649 144351 331726
rect 121706 16020 124408 331649
rect 147278 329206 149690 366112
rect 121706 15580 122810 16020
rect 123250 15580 124408 16020
rect 121706 15520 124408 15580
rect 121706 15080 122810 15520
rect 123250 15080 124408 15520
rect 121706 15020 124408 15080
rect 121706 14580 122810 15020
rect 123250 14580 124408 15020
rect 121706 14520 124408 14580
rect 121706 14080 122810 14520
rect 123250 14080 124408 14520
rect 121706 14020 124408 14080
rect 121706 13580 122810 14020
rect 123250 13580 124408 14020
rect 121706 13520 124408 13580
rect 121706 13080 122810 13520
rect 123250 13080 124408 13520
rect 121706 13020 124408 13080
rect 121706 12580 122810 13020
rect 123250 12580 124408 13020
rect 121706 12520 124408 12580
rect 121706 12080 122810 12520
rect 123250 12080 124408 12520
rect 121706 12000 124408 12080
rect 126266 326794 149690 329206
rect 126266 16020 128678 326794
rect 151416 324430 154276 363246
rect 126266 15580 127240 16020
rect 127680 15580 128678 16020
rect 126266 15520 128678 15580
rect 126266 15080 127240 15520
rect 127680 15080 128678 15520
rect 126266 15020 128678 15080
rect 126266 14580 127240 15020
rect 127680 14580 128678 15020
rect 126266 14520 128678 14580
rect 126266 14080 127240 14520
rect 127680 14080 128678 14520
rect 126266 14020 128678 14080
rect 126266 13580 127240 14020
rect 127680 13580 128678 14020
rect 126266 13520 128678 13580
rect 126266 13080 127240 13520
rect 127680 13080 128678 13520
rect 126266 13020 128678 13080
rect 126266 12580 127240 13020
rect 127680 12580 128678 13020
rect 126266 12520 128678 12580
rect 126266 12080 127240 12520
rect 127680 12080 128678 12520
rect 126266 12000 128678 12080
rect 130404 321570 154276 324430
rect 130404 16020 133264 321570
rect 155944 319368 158680 359426
rect 130404 15580 131600 16020
rect 132040 15580 133264 16020
rect 130404 15520 133264 15580
rect 130404 15080 131600 15520
rect 132040 15080 133264 15520
rect 130404 15020 133264 15080
rect 130404 14580 131600 15020
rect 132040 14580 133264 15020
rect 130404 14520 133264 14580
rect 130404 14080 131600 14520
rect 132040 14080 133264 14520
rect 130404 14020 133264 14080
rect 130404 13580 131600 14020
rect 132040 13580 133264 14020
rect 130404 13520 133264 13580
rect 130404 13080 131600 13520
rect 132040 13080 133264 13520
rect 130404 13020 133264 13080
rect 130404 12580 131600 13020
rect 132040 12580 133264 13020
rect 130404 12520 133264 12580
rect 130404 12080 131600 12520
rect 132040 12080 133264 12520
rect 130404 12000 133264 12080
rect 134932 316632 158680 319368
rect 134932 16020 137668 316632
rect 160188 313000 163156 356244
rect 139176 310032 163156 313000
rect 139176 35150 142144 310032
rect 164902 307000 167546 352407
rect 185904 315880 188762 329656
rect 185904 315580 185912 315880
rect 186212 315580 186272 315880
rect 186572 315580 186632 315880
rect 186932 315580 186992 315880
rect 187292 315580 187352 315880
rect 187652 315580 187712 315880
rect 188012 315580 188072 315880
rect 188372 315580 188432 315880
rect 188732 315580 188762 315880
rect 185904 315520 188762 315580
rect 185904 315220 185912 315520
rect 186212 315220 186272 315520
rect 186572 315220 186632 315520
rect 186932 315220 186992 315520
rect 187292 315220 187352 315520
rect 187652 315220 187712 315520
rect 188012 315220 188072 315520
rect 188372 315220 188432 315520
rect 188732 315220 188762 315520
rect 185904 315160 188762 315220
rect 185904 314860 185912 315160
rect 186212 314860 186272 315160
rect 186572 314860 186632 315160
rect 186932 314860 186992 315160
rect 187292 314860 187352 315160
rect 187652 314860 187712 315160
rect 188012 314860 188072 315160
rect 188372 314860 188432 315160
rect 188732 314860 188762 315160
rect 185904 314800 188762 314860
rect 185904 314500 185912 314800
rect 186212 314500 186272 314800
rect 186572 314500 186632 314800
rect 186932 314500 186992 314800
rect 187292 314500 187352 314800
rect 187652 314500 187712 314800
rect 188012 314500 188072 314800
rect 188372 314500 188432 314800
rect 188732 314500 188762 314800
rect 185904 314440 188762 314500
rect 185904 314140 185912 314440
rect 186212 314140 186272 314440
rect 186572 314140 186632 314440
rect 186932 314140 186992 314440
rect 187292 314140 187352 314440
rect 187652 314140 187712 314440
rect 188012 314140 188072 314440
rect 188372 314140 188432 314440
rect 188732 314140 188762 314440
rect 185904 314080 188762 314140
rect 185904 313780 185912 314080
rect 186212 313780 186272 314080
rect 186572 313780 186632 314080
rect 186932 313780 186992 314080
rect 187292 313780 187352 314080
rect 187652 313780 187712 314080
rect 188012 313780 188072 314080
rect 188372 313780 188432 314080
rect 188732 313780 188762 314080
rect 185904 313760 188762 313780
rect 261726 310414 264584 328411
rect 261726 310114 261734 310414
rect 262034 310114 262094 310414
rect 262394 310114 262454 310414
rect 262754 310114 262814 310414
rect 263114 310114 263174 310414
rect 263474 310114 263534 310414
rect 263834 310114 263894 310414
rect 264194 310114 264254 310414
rect 264554 310114 264584 310414
rect 261726 310054 264584 310114
rect 261726 309754 261734 310054
rect 262034 309754 262094 310054
rect 262394 309754 262454 310054
rect 262754 309754 262814 310054
rect 263114 309754 263174 310054
rect 263474 309754 263534 310054
rect 263834 309754 263894 310054
rect 264194 309754 264254 310054
rect 264554 309754 264584 310054
rect 261726 309694 264584 309754
rect 261726 309394 261734 309694
rect 262034 309394 262094 309694
rect 262394 309394 262454 309694
rect 262754 309394 262814 309694
rect 263114 309394 263174 309694
rect 263474 309394 263534 309694
rect 263834 309394 263894 309694
rect 264194 309394 264254 309694
rect 264554 309394 264584 309694
rect 261726 309334 264584 309394
rect 261726 309034 261734 309334
rect 262034 309034 262094 309334
rect 262394 309034 262454 309334
rect 262754 309034 262814 309334
rect 263114 309034 263174 309334
rect 263474 309034 263534 309334
rect 263834 309034 263894 309334
rect 264194 309034 264254 309334
rect 264554 309034 264584 309334
rect 261726 308974 264584 309034
rect 261726 308674 261734 308974
rect 262034 308674 262094 308974
rect 262394 308674 262454 308974
rect 262754 308674 262814 308974
rect 263114 308674 263174 308974
rect 263474 308674 263534 308974
rect 263834 308674 263894 308974
rect 264194 308674 264254 308974
rect 264554 308674 264584 308974
rect 261726 308614 264584 308674
rect 261726 308314 261734 308614
rect 262034 308314 262094 308614
rect 262394 308314 262454 308614
rect 262754 308314 262814 308614
rect 263114 308314 263174 308614
rect 263474 308314 263534 308614
rect 263834 308314 263894 308614
rect 264194 308314 264254 308614
rect 264554 308314 264584 308614
rect 261726 308280 264584 308314
rect 139176 34550 139200 35150
rect 139800 34550 139960 35150
rect 140560 34550 140740 35150
rect 141340 34550 141500 35150
rect 142100 34550 142144 35150
rect 139176 34450 142144 34550
rect 143472 304356 167546 307000
rect 134932 15580 136080 16020
rect 136520 15580 137668 16020
rect 134932 15520 137668 15580
rect 134932 15080 136080 15520
rect 136520 15080 137668 15520
rect 134932 15020 137668 15080
rect 134932 14580 136080 15020
rect 136520 14580 137668 15020
rect 134932 14520 137668 14580
rect 134932 14080 136080 14520
rect 136520 14080 137668 14520
rect 134932 14020 137668 14080
rect 134932 13580 136080 14020
rect 136520 13580 137668 14020
rect 134932 13520 137668 13580
rect 134932 13080 136080 13520
rect 136520 13080 137668 13520
rect 134932 13020 137668 13080
rect 134932 12580 136080 13020
rect 136520 12580 137668 13020
rect 134932 12520 137668 12580
rect 134932 12080 136080 12520
rect 136520 12080 137668 12520
rect 134932 12000 137668 12080
rect 143472 14520 146116 304356
rect 339520 304188 342378 332534
rect 339520 303888 339528 304188
rect 339828 303888 339888 304188
rect 340188 303888 340248 304188
rect 340548 303888 340608 304188
rect 340908 303888 340968 304188
rect 341268 303888 341328 304188
rect 341628 303888 341688 304188
rect 341988 303888 342048 304188
rect 342348 303888 342378 304188
rect 339520 303828 342378 303888
rect 339520 303528 339528 303828
rect 339828 303528 339888 303828
rect 340188 303528 340248 303828
rect 340548 303528 340608 303828
rect 340908 303528 340968 303828
rect 341268 303528 341328 303828
rect 341628 303528 341688 303828
rect 341988 303528 342048 303828
rect 342348 303528 342378 303828
rect 339520 303468 342378 303528
rect 339520 303168 339528 303468
rect 339828 303168 339888 303468
rect 340188 303168 340248 303468
rect 340548 303168 340608 303468
rect 340908 303168 340968 303468
rect 341268 303168 341328 303468
rect 341628 303168 341688 303468
rect 341988 303168 342048 303468
rect 342348 303168 342378 303468
rect 339520 303108 342378 303168
rect 339520 302808 339528 303108
rect 339828 302808 339888 303108
rect 340188 302808 340248 303108
rect 340548 302808 340608 303108
rect 340908 302808 340968 303108
rect 341268 302808 341328 303108
rect 341628 302808 341688 303108
rect 341988 302808 342048 303108
rect 342348 302808 342378 303108
rect 339520 302748 342378 302808
rect 339520 302448 339528 302748
rect 339828 302448 339888 302748
rect 340188 302448 340248 302748
rect 340548 302448 340608 302748
rect 340908 302448 340968 302748
rect 341268 302448 341328 302748
rect 341628 302448 341688 302748
rect 341988 302448 342048 302748
rect 342348 302448 342378 302748
rect 339520 302388 342378 302448
rect 339520 302088 339528 302388
rect 339828 302088 339888 302388
rect 340188 302088 340248 302388
rect 340548 302088 340608 302388
rect 340908 302088 340968 302388
rect 341268 302088 341328 302388
rect 341628 302088 341688 302388
rect 341988 302088 342048 302388
rect 342348 302088 342378 302388
rect 339520 302020 342378 302088
rect 542000 47401 543000 486200
rect 544000 361980 545000 488000
rect 544001 92201 545000 361980
rect 546000 272201 547000 490000
rect 548000 316601 549000 492200
rect 550000 359801 552000 568999
rect 553000 405601 553400 572999
rect 555000 450001 555400 574999
rect 568000 500400 574000 589200
rect 568000 499800 568200 500400
rect 568800 499800 569000 500400
rect 569600 499800 569800 500400
rect 570400 499800 570600 500400
rect 571200 499800 571400 500400
rect 572000 499800 572200 500400
rect 572800 499800 573000 500400
rect 573600 499800 574000 500400
rect 568000 456000 574000 499800
rect 568000 455400 568200 456000
rect 568800 455400 569000 456000
rect 569600 455400 569800 456000
rect 570400 455400 570600 456000
rect 571200 455400 571400 456000
rect 572000 455400 572200 456000
rect 572800 455400 573000 456000
rect 573600 455400 574000 456000
rect 554999 450000 555401 450001
rect 554999 449600 555000 450000
rect 555400 449600 555401 450000
rect 554999 449599 555401 449600
rect 568000 411600 574000 455400
rect 568000 411000 568200 411600
rect 568800 411000 569000 411600
rect 569600 411000 569800 411600
rect 570400 411000 570600 411600
rect 571200 411000 571400 411600
rect 572000 411000 572200 411600
rect 572800 411000 573000 411600
rect 573600 411000 574000 411600
rect 552999 405600 553401 405601
rect 552999 405200 553000 405600
rect 553400 405200 553401 405600
rect 552999 405199 553401 405200
rect 568000 365200 574000 411000
rect 568000 364600 568200 365200
rect 568800 364600 569000 365200
rect 569600 364600 569800 365200
rect 570400 364600 570600 365200
rect 571200 364600 571400 365200
rect 572000 364600 572200 365200
rect 572800 364600 573000 365200
rect 573600 364600 574000 365200
rect 568000 364400 574000 364600
rect 549999 359800 552001 359801
rect 549999 357800 550000 359800
rect 552000 357800 552001 359800
rect 549999 357799 552001 357800
rect 547999 316600 549001 316601
rect 547999 315600 548000 316600
rect 549000 315600 549001 316600
rect 547999 315599 549001 315600
rect 545999 272200 547001 272201
rect 545999 271200 546000 272200
rect 547000 271200 547001 272200
rect 545999 271199 547001 271200
rect 543999 92200 545001 92201
rect 543999 91200 544000 92200
rect 545000 91200 545001 92200
rect 543999 91199 545001 91200
rect 541999 47400 543001 47401
rect 541999 46400 542000 47400
rect 543000 46400 543001 47400
rect 541999 46399 543001 46400
rect 143472 14080 144562 14520
rect 145002 14080 146116 14520
rect 143472 14020 146116 14080
rect 143472 13580 144562 14020
rect 145002 13580 146116 14020
rect 143472 13520 146116 13580
rect 143472 13080 144562 13520
rect 145002 13080 146116 13520
rect 143472 13020 146116 13080
rect 143472 12580 144562 13020
rect 145002 12580 146116 13020
rect 143472 12520 146116 12580
rect 143472 12080 144562 12520
rect 145002 12080 146116 12520
rect 143472 12000 146116 12080
<< rmetal4 >>
rect 524200 677300 528400 679300
rect 35000 181000 41000 197114
<< via4 >>
rect 177000 698800 179400 699000
rect 177000 696800 177200 698800
rect 177200 696800 179200 698800
rect 179200 696800 179400 698800
rect 177000 696600 179400 696800
rect 228600 698900 231000 699000
rect 228600 696700 228700 698900
rect 228700 696700 230900 698900
rect 230900 696700 231000 698900
rect 228600 696600 231000 696700
rect 7600 567200 12400 567400
rect 7600 563800 7800 567200
rect 7800 563800 12200 567200
rect 12200 563800 12400 567200
rect 7600 563600 12400 563800
rect 7600 563000 12400 563200
rect 7600 559600 7800 563000
rect 7800 559600 12200 563000
rect 12200 559600 12400 563000
rect 7600 559400 12400 559600
rect 389600 559600 397400 567200
rect 20200 521200 27800 528800
rect 10000 505200 11000 506200
rect 11200 505200 12200 506200
rect 12400 505200 13400 506200
rect 13600 505200 14600 506200
rect 14800 505200 15800 506200
rect 34200 504200 41800 511800
rect 10000 462000 11000 463000
rect 11200 462000 12200 463000
rect 12400 462000 13400 463000
rect 13600 462000 14600 463000
rect 14800 462000 15800 463000
rect 10000 418800 11000 419800
rect 11200 418800 12200 419800
rect 12400 418800 13400 419800
rect 13600 418800 14600 419800
rect 14800 418800 15800 419800
rect 10000 375400 11000 376400
rect 11200 375400 12200 376400
rect 12400 375400 13400 376400
rect 13600 375400 14600 376400
rect 14800 375400 15800 376400
rect 10000 332200 11000 333200
rect 11200 332200 12200 333200
rect 12400 332200 13400 333200
rect 13600 332200 14600 333200
rect 14800 332200 15800 333200
rect 10000 289000 11000 290000
rect 11200 289000 12200 290000
rect 12400 289000 13400 290000
rect 13600 289000 14600 290000
rect 14800 289000 15800 290000
rect 10000 246000 11000 247000
rect 11200 246000 12200 247000
rect 12400 246000 13400 247000
rect 13600 246000 14600 247000
rect 14800 246000 15800 247000
rect 117500 369100 120100 370900
rect 60080 346300 60680 346310
rect 60080 345740 60100 346300
rect 60100 345740 60660 346300
rect 60660 345740 60680 346300
rect 60080 345710 60680 345740
rect 60780 346300 61380 346310
rect 60780 345740 60800 346300
rect 60800 345740 61360 346300
rect 61360 345740 61380 346300
rect 60780 345710 61380 345740
rect 61480 346300 62080 346310
rect 61480 345740 61500 346300
rect 61500 345740 62060 346300
rect 62060 345740 62080 346300
rect 61480 345710 62080 345740
rect 62180 346300 62780 346310
rect 62180 345740 62200 346300
rect 62200 345740 62760 346300
rect 62760 345740 62780 346300
rect 62180 345710 62780 345740
rect 60080 345600 60680 345610
rect 60080 345040 60100 345600
rect 60100 345040 60660 345600
rect 60660 345040 60680 345600
rect 60080 345010 60680 345040
rect 60780 345600 61380 345610
rect 60780 345040 60800 345600
rect 60800 345040 61360 345600
rect 61360 345040 61380 345600
rect 60780 345010 61380 345040
rect 61480 345600 62080 345610
rect 61480 345040 61500 345600
rect 61500 345040 62060 345600
rect 62060 345040 62080 345600
rect 61480 345010 62080 345040
rect 62180 345600 62780 345610
rect 62180 345040 62200 345600
rect 62200 345040 62760 345600
rect 62760 345040 62780 345600
rect 62180 345010 62780 345040
rect 60080 344900 60680 344910
rect 60080 344340 60100 344900
rect 60100 344340 60660 344900
rect 60660 344340 60680 344900
rect 60080 344310 60680 344340
rect 60780 344900 61380 344910
rect 60780 344340 60800 344900
rect 60800 344340 61360 344900
rect 61360 344340 61380 344900
rect 60780 344310 61380 344340
rect 61480 344900 62080 344910
rect 61480 344340 61500 344900
rect 61500 344340 62060 344900
rect 62060 344340 62080 344900
rect 61480 344310 62080 344340
rect 62180 344900 62780 344910
rect 62180 344340 62200 344900
rect 62200 344340 62760 344900
rect 62760 344340 62780 344900
rect 62180 344310 62780 344340
rect 60052 342814 60652 342824
rect 60052 342254 60072 342814
rect 60072 342254 60632 342814
rect 60632 342254 60652 342814
rect 60052 342224 60652 342254
rect 60752 342814 61352 342824
rect 60752 342254 60772 342814
rect 60772 342254 61332 342814
rect 61332 342254 61352 342814
rect 60752 342224 61352 342254
rect 61452 342814 62052 342824
rect 61452 342254 61472 342814
rect 61472 342254 62032 342814
rect 62032 342254 62052 342814
rect 61452 342224 62052 342254
rect 62152 342814 62752 342824
rect 62152 342254 62172 342814
rect 62172 342254 62732 342814
rect 62732 342254 62752 342814
rect 62152 342224 62752 342254
rect 60052 342114 60652 342124
rect 60052 341554 60072 342114
rect 60072 341554 60632 342114
rect 60632 341554 60652 342114
rect 60052 341524 60652 341554
rect 60752 342114 61352 342124
rect 60752 341554 60772 342114
rect 60772 341554 61332 342114
rect 61332 341554 61352 342114
rect 60752 341524 61352 341554
rect 61452 342114 62052 342124
rect 61452 341554 61472 342114
rect 61472 341554 62032 342114
rect 62032 341554 62052 342114
rect 61452 341524 62052 341554
rect 62152 342114 62752 342124
rect 62152 341554 62172 342114
rect 62172 341554 62732 342114
rect 62732 341554 62752 342114
rect 62152 341524 62752 341554
rect 60052 341414 60652 341424
rect 60052 340854 60072 341414
rect 60072 340854 60632 341414
rect 60632 340854 60652 341414
rect 60052 340824 60652 340854
rect 60752 341414 61352 341424
rect 60752 340854 60772 341414
rect 60772 340854 61332 341414
rect 61332 340854 61352 341414
rect 60752 340824 61352 340854
rect 61452 341414 62052 341424
rect 61452 340854 61472 341414
rect 61472 340854 62032 341414
rect 62032 340854 62052 341414
rect 61452 340824 62052 340854
rect 62152 341414 62752 341424
rect 62152 340854 62172 341414
rect 62172 340854 62732 341414
rect 62732 340854 62752 341414
rect 62152 340824 62752 340854
rect 60120 339174 60720 339184
rect 60120 338614 60140 339174
rect 60140 338614 60700 339174
rect 60700 338614 60720 339174
rect 60120 338584 60720 338614
rect 60820 339174 61420 339184
rect 60820 338614 60840 339174
rect 60840 338614 61400 339174
rect 61400 338614 61420 339174
rect 60820 338584 61420 338614
rect 61520 339174 62120 339184
rect 61520 338614 61540 339174
rect 61540 338614 62100 339174
rect 62100 338614 62120 339174
rect 61520 338584 62120 338614
rect 62220 339174 62820 339184
rect 62220 338614 62240 339174
rect 62240 338614 62800 339174
rect 62800 338614 62820 339174
rect 62220 338584 62820 338614
rect 60120 338474 60720 338484
rect 60120 337914 60140 338474
rect 60140 337914 60700 338474
rect 60700 337914 60720 338474
rect 60120 337884 60720 337914
rect 60820 338474 61420 338484
rect 60820 337914 60840 338474
rect 60840 337914 61400 338474
rect 61400 337914 61420 338474
rect 60820 337884 61420 337914
rect 61520 338474 62120 338484
rect 61520 337914 61540 338474
rect 61540 337914 62100 338474
rect 62100 337914 62120 338474
rect 61520 337884 62120 337914
rect 62220 338474 62820 338484
rect 62220 337914 62240 338474
rect 62240 337914 62800 338474
rect 62800 337914 62820 338474
rect 62220 337884 62820 337914
rect 60120 337774 60720 337784
rect 60120 337214 60140 337774
rect 60140 337214 60700 337774
rect 60700 337214 60720 337774
rect 60120 337184 60720 337214
rect 60820 337774 61420 337784
rect 60820 337214 60840 337774
rect 60840 337214 61400 337774
rect 61400 337214 61420 337774
rect 60820 337184 61420 337214
rect 61520 337774 62120 337784
rect 61520 337214 61540 337774
rect 61540 337214 62100 337774
rect 62100 337214 62120 337774
rect 61520 337184 62120 337214
rect 62220 337774 62820 337784
rect 62220 337214 62240 337774
rect 62240 337214 62800 337774
rect 62800 337214 62820 337774
rect 62220 337184 62820 337214
rect 60120 335070 60720 335080
rect 60120 334510 60140 335070
rect 60140 334510 60700 335070
rect 60700 334510 60720 335070
rect 60120 334480 60720 334510
rect 60820 335070 61420 335080
rect 60820 334510 60840 335070
rect 60840 334510 61400 335070
rect 61400 334510 61420 335070
rect 60820 334480 61420 334510
rect 61520 335070 62120 335080
rect 61520 334510 61540 335070
rect 61540 334510 62100 335070
rect 62100 334510 62120 335070
rect 61520 334480 62120 334510
rect 62220 335070 62820 335080
rect 62220 334510 62240 335070
rect 62240 334510 62800 335070
rect 62800 334510 62820 335070
rect 62220 334480 62820 334510
rect 60120 334370 60720 334380
rect 60120 333810 60140 334370
rect 60140 333810 60700 334370
rect 60700 333810 60720 334370
rect 60120 333780 60720 333810
rect 60820 334370 61420 334380
rect 60820 333810 60840 334370
rect 60840 333810 61400 334370
rect 61400 333810 61420 334370
rect 60820 333780 61420 333810
rect 61520 334370 62120 334380
rect 61520 333810 61540 334370
rect 61540 333810 62100 334370
rect 62100 333810 62120 334370
rect 61520 333780 62120 333810
rect 62220 334370 62820 334380
rect 62220 333810 62240 334370
rect 62240 333810 62800 334370
rect 62800 333810 62820 334370
rect 62220 333780 62820 333810
rect 60120 333670 60720 333680
rect 60120 333110 60140 333670
rect 60140 333110 60700 333670
rect 60700 333110 60720 333670
rect 60120 333080 60720 333110
rect 60820 333670 61420 333680
rect 60820 333110 60840 333670
rect 60840 333110 61400 333670
rect 61400 333110 61420 333670
rect 60820 333080 61420 333110
rect 61520 333670 62120 333680
rect 61520 333110 61540 333670
rect 61540 333110 62100 333670
rect 62100 333110 62120 333670
rect 61520 333080 62120 333110
rect 62220 333670 62820 333680
rect 62220 333110 62240 333670
rect 62240 333110 62800 333670
rect 62800 333110 62820 333670
rect 62220 333080 62820 333110
rect 60120 331624 60720 331634
rect 60120 331064 60140 331624
rect 60140 331064 60700 331624
rect 60700 331064 60720 331624
rect 60120 331034 60720 331064
rect 60820 331624 61420 331634
rect 60820 331064 60840 331624
rect 60840 331064 61400 331624
rect 61400 331064 61420 331624
rect 60820 331034 61420 331064
rect 61520 331624 62120 331634
rect 61520 331064 61540 331624
rect 61540 331064 62100 331624
rect 62100 331064 62120 331624
rect 61520 331034 62120 331064
rect 62220 331624 62820 331634
rect 62220 331064 62240 331624
rect 62240 331064 62800 331624
rect 62800 331064 62820 331624
rect 62220 331034 62820 331064
rect 60120 330924 60720 330934
rect 60120 330364 60140 330924
rect 60140 330364 60700 330924
rect 60700 330364 60720 330924
rect 60120 330334 60720 330364
rect 60820 330924 61420 330934
rect 60820 330364 60840 330924
rect 60840 330364 61400 330924
rect 61400 330364 61420 330924
rect 60820 330334 61420 330364
rect 61520 330924 62120 330934
rect 61520 330364 61540 330924
rect 61540 330364 62100 330924
rect 62100 330364 62120 330924
rect 61520 330334 62120 330364
rect 62220 330924 62820 330934
rect 62220 330364 62240 330924
rect 62240 330364 62800 330924
rect 62800 330364 62820 330924
rect 62220 330334 62820 330364
rect 60120 330224 60720 330234
rect 60120 329664 60140 330224
rect 60140 329664 60700 330224
rect 60700 329664 60720 330224
rect 60120 329634 60720 329664
rect 60820 330224 61420 330234
rect 60820 329664 60840 330224
rect 60840 329664 61400 330224
rect 61400 329664 61420 330224
rect 60820 329634 61420 329664
rect 61520 330224 62120 330234
rect 61520 329664 61540 330224
rect 61540 329664 62100 330224
rect 62100 329664 62120 330224
rect 61520 329634 62120 329664
rect 62220 330224 62820 330234
rect 62220 329664 62240 330224
rect 62240 329664 62800 330224
rect 62800 329664 62820 330224
rect 62220 329634 62820 329664
rect 10000 118400 11000 119400
rect 11200 118400 12200 119400
rect 12400 118400 13400 119400
rect 13600 118400 14600 119400
rect 14800 118400 15800 119400
rect 10000 75200 11000 76200
rect 11200 75200 12200 76200
rect 12400 75200 13400 76200
rect 13600 75200 14600 76200
rect 14800 75200 15800 76200
<< metal5 >>
rect 165594 700000 170594 704800
rect 175894 700000 180894 704800
rect 165594 699000 180894 700000
rect 165594 696600 177000 699000
rect 179400 696600 180894 699000
rect 165594 695150 180894 696600
rect 217294 700000 222294 704800
rect 227594 700000 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 217294 699000 232594 700000
rect 217294 696600 228600 699000
rect 231000 696600 232594 699000
rect 169200 642000 177200 695150
rect 217294 695100 232594 696600
rect 221000 654000 229000 695100
rect 221000 646000 438400 654000
rect 169200 634000 430000 642000
rect 430400 625692 438400 646000
rect 7576 567400 12424 567424
rect 7400 563600 7600 567400
rect 12400 563600 16400 567400
rect 7400 563200 16400 563600
rect 7400 559400 7600 563200
rect 12400 559400 16400 563200
rect 20400 567200 397623 567400
rect 20400 559600 389600 567200
rect 397400 559600 397623 567200
rect 20400 559400 397623 559600
rect 7576 559376 12424 559400
rect 20000 528800 28000 529000
rect 20000 528000 20200 528800
rect 10000 522000 20200 528000
rect 10001 506224 16000 522000
rect 20000 521200 20200 522000
rect 27800 528000 28000 528800
rect 27800 522000 52000 528000
rect 27800 521200 28000 522000
rect 20000 521000 28000 521200
rect 9976 506200 16000 506224
rect 9976 505200 10000 506200
rect 11000 505200 11200 506200
rect 12200 505200 12400 506200
rect 13400 505200 13600 506200
rect 14600 505200 14800 506200
rect 15800 505200 16000 506200
rect 9976 505176 16000 505200
rect 10001 463024 16000 505176
rect 34000 511800 53000 512000
rect 34000 504200 34200 511800
rect 41800 504200 53000 511800
rect 34000 504000 53000 504200
rect 9976 463000 16000 463024
rect 9976 462000 10000 463000
rect 11000 462000 11200 463000
rect 12200 462000 12400 463000
rect 13400 462000 13600 463000
rect 14600 462000 14800 463000
rect 15800 462000 16000 463000
rect 9976 461976 16000 462000
rect 10001 419824 16000 461976
rect 9976 419800 16000 419824
rect 9976 418800 10000 419800
rect 11000 418800 11200 419800
rect 12200 418800 12400 419800
rect 13400 418800 13600 419800
rect 14600 418800 14800 419800
rect 15800 418800 16000 419800
rect 9976 418776 16000 418800
rect 10001 376424 16000 418776
rect 9976 376400 16000 376424
rect 9976 375400 10000 376400
rect 11000 375400 11200 376400
rect 12200 375400 12400 376400
rect 13400 375400 13600 376400
rect 14600 375400 14800 376400
rect 15800 375400 16000 376400
rect 9976 375376 16000 375400
rect 10001 333224 16000 375376
rect 117476 370900 120124 370924
rect 117476 369100 117500 370900
rect 120100 369100 120124 370900
rect 117476 369076 120124 369100
rect 60040 346310 62820 346350
rect 60040 345710 60080 346310
rect 60680 345710 60780 346310
rect 61380 345710 61480 346310
rect 62080 345710 62180 346310
rect 62780 345710 62820 346310
rect 60040 345610 62820 345710
rect 60040 345010 60080 345610
rect 60680 345010 60780 345610
rect 61380 345010 61480 345610
rect 62080 345010 62180 345610
rect 62780 345010 62820 345610
rect 60040 344910 62820 345010
rect 60040 344310 60080 344910
rect 60680 344310 60780 344910
rect 61380 344310 61480 344910
rect 62080 344310 62180 344910
rect 62780 344310 62820 344910
rect 60040 344280 62820 344310
rect 60012 342824 62792 342864
rect 60012 342224 60052 342824
rect 60652 342224 60752 342824
rect 61352 342224 61452 342824
rect 62052 342224 62152 342824
rect 62752 342224 62792 342824
rect 60012 342124 62792 342224
rect 60012 341524 60052 342124
rect 60652 341524 60752 342124
rect 61352 341524 61452 342124
rect 62052 341524 62152 342124
rect 62752 341524 62792 342124
rect 60012 341424 62792 341524
rect 60012 340824 60052 341424
rect 60652 340824 60752 341424
rect 61352 340824 61452 341424
rect 62052 340824 62152 341424
rect 62752 340824 62792 341424
rect 60012 340794 62792 340824
rect 60080 339184 62860 339224
rect 60080 338584 60120 339184
rect 60720 338584 60820 339184
rect 61420 338584 61520 339184
rect 62120 338584 62220 339184
rect 62820 338584 62860 339184
rect 60080 338484 62860 338584
rect 60080 337884 60120 338484
rect 60720 337884 60820 338484
rect 61420 337884 61520 338484
rect 62120 337884 62220 338484
rect 62820 337884 62860 338484
rect 60080 337784 62860 337884
rect 60080 337184 60120 337784
rect 60720 337184 60820 337784
rect 61420 337184 61520 337784
rect 62120 337184 62220 337784
rect 62820 337184 62860 337784
rect 60080 337154 62860 337184
rect 9976 333200 16000 333224
rect 9976 332200 10000 333200
rect 11000 332200 11200 333200
rect 12200 332200 12400 333200
rect 13400 332200 13600 333200
rect 14600 332200 14800 333200
rect 15800 332200 16000 333200
rect 60080 335080 62860 335120
rect 60080 334480 60120 335080
rect 60720 334480 60820 335080
rect 61420 334480 61520 335080
rect 62120 334480 62220 335080
rect 62820 334480 62860 335080
rect 60080 334380 62860 334480
rect 60080 333780 60120 334380
rect 60720 333780 60820 334380
rect 61420 333780 61520 334380
rect 62120 333780 62220 334380
rect 62820 333780 62860 334380
rect 60080 333680 62860 333780
rect 60080 333080 60120 333680
rect 60720 333080 60820 333680
rect 61420 333080 61520 333680
rect 62120 333080 62220 333680
rect 62820 333080 62860 333680
rect 60080 333050 62860 333080
rect 9976 332176 16000 332200
rect 10001 290024 16000 332176
rect 60080 331634 62860 331674
rect 60080 331034 60120 331634
rect 60720 331034 60820 331634
rect 61420 331034 61520 331634
rect 62120 331034 62220 331634
rect 62820 331034 62860 331634
rect 60080 330934 62860 331034
rect 60080 330334 60120 330934
rect 60720 330334 60820 330934
rect 61420 330334 61520 330934
rect 62120 330334 62220 330934
rect 62820 330334 62860 330934
rect 60080 330234 62860 330334
rect 60080 329634 60120 330234
rect 60720 329634 60820 330234
rect 61420 329634 61520 330234
rect 62120 329634 62220 330234
rect 62820 329634 62860 330234
rect 60080 329604 62860 329634
rect 9976 290000 16000 290024
rect 9976 289000 10000 290000
rect 11000 289000 11200 290000
rect 12200 289000 12400 290000
rect 13400 289000 13600 290000
rect 14600 289000 14800 290000
rect 15800 289000 16000 290000
rect 9976 288976 16000 289000
rect 10001 247024 16000 288976
rect 9976 247000 16000 247024
rect 9976 246000 10000 247000
rect 11000 246000 11200 247000
rect 12200 246000 12400 247000
rect 13400 246000 13600 247000
rect 14600 246000 14800 247000
rect 15800 246000 16000 247000
rect 9976 245976 16000 246000
rect 10001 119424 16000 245976
rect 9976 119400 16000 119424
rect 9976 118400 10000 119400
rect 11000 118400 11200 119400
rect 12200 118400 12400 119400
rect 13400 118400 13600 119400
rect 14600 118400 14800 119400
rect 15800 118400 16000 119400
rect 9976 118376 16000 118400
rect 10001 76224 16000 118376
rect 9976 76200 16000 76224
rect 9976 75200 10000 76200
rect 11000 75200 11200 76200
rect 12200 75200 12400 76200
rect 13400 75200 13600 76200
rect 14600 75200 14800 76200
rect 15800 75200 16000 76200
rect 9976 75176 16000 75200
rect 10001 75100 16000 75176
<< rm5 >>
rect 16400 559400 20400 567400
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 49000 654000 535000 655000
rect 49000 50000 50000 654000
rect 534000 50000 535000 654000
rect 49000 49000 535000 50000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use dac_top_cell  dac_top_cell_0 ../user_prj/UNIC-CASS_precheck_dac/mag
timestamp 1699094506
transform 1 0 503758 0 1 525566
box -28028 -20682 27930 18344
use MulColROs  MulColROs_0 ../user_prj/MulColRO/mag
timestamp 1699009326
transform 1 0 -11386 0 1 -273116
box 62168 599934 367990 811050
use ulqc_ldo  ulqc_ldo_0 ../user_prj/ULQC_LDO/mag
timestamp 1699276451
transform 1 0 387749 0 1 602932
box -2065 -11200 50651 31068
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
